XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��)�t�@�*������N�	��h����
p\���~�(r�!��p![����puj��@{g�d9���u��@o�	���\��j�{��b���@�gq5��O�o*�'�-Ӳ��[��d����$��к�UJ�%��SgY~�:�A|<�ӣS�}�%�C�n0��f�7��S3�Ї��_�F�1m  �]^T
�8��;��#A�i!Z���\l�%D0f����aiHQ�4ěőG�5�/�.ÈP�]=��&ӆ����G!����ט�F,��_�ׯc�W��n�	ŕpv�Ҥ|5��%����C� ���$2$�k�>3o��infrb8�P�E�rM�8�"�Jxl����C��I	nRf�Y���81��Ǥ��r;���];�\h��dMX&B9��<��QD���u�X�B?V�ozv͵�fz*�v�հ���^6�\�e�*�U(u��[i��\33���}���M��|��C�&#��u����| ��uP|W��y�"���&�8Ķ#������sn�b�,�NT�ߎ:�My[A��Pi)�~���yh�ˋ��*(�Z�M���bC}C�`�k��	��\ �C?.z�d&��D��,�.Q5u~8&i_�*y�M�.�ѷ���ma��=��T��,��8+rB~��6	�I����-��9��JdA��H4��j�R�U �Qr��p��T��!���<� ����gʽ�IfO��7AזA����Kx1�i(2u[�ی`%��O�����:���.XlxVHYEB    3fdc    1160���p1�ܕT2��'��̘l���l�"�>��.��TD��nx�y=l&�خ�Ei e8-|�Zw4~�mT)��+x1�L�m�zj[4�>&�Iv��r(��=���HcTmB*��r���gE��x'�Թ�^ 	�S_��׍���zk]$�)�I�W�*D�{o�q�Q���Ai� ���_
�U�Q���.=����| �c6]ܷ���WH��C+�E�w>}�v/�c��\;���y���&:�6Ko7Ro�i��ѶT��U�^�!.���@� 
@���i۝��!����x67��v�����[�0�Tä�7�N�!�^��E�I����#tgM��ϓW�fH�Aq�#ZǴw�V-��>�����+����OZ�n�]���&���[9��1SBH������b�Eo���[r��Jq�����@�K�bR�'������Y��Zw�����#���S�q�KiD(��IA|�J��&ʊ�Y�_�wt$��mY�ByϨ�7ff`�7&̼nqu٦�v3H�9Wn޹�^hr�a����o%��;�X���5Nޅ'����e��֋+�[��<.E�(�� 1��XA�:��c�?d�A���E��|G��vsk��!�R4	�5N @���!B����Ȏ�f�����u��O�/�x���dl~A���	�`
Y���M|/����Ǭ~�#�p��j��MѦ��ZZw�Ze?aJ��?���yoX��L�U��9��zp�-3�Vn,�]㫐Q�F�X}����Z���.9�7C\Xii����O���%�/.,r�2�R6��u�~h��ĒX�Bd������B �����/��[:�$� ��;!��'d���G�C�-z~/��Z\�D9���y��+���77����:��Ԧ��3�7����"u���S�p��L���H�e�6�?w@Z�֐	�\�ǔC�(!���Q� ����n��b{�_)����ë�)��#�����c P )��X������H�{�NU�C��
�f	o�.l��V��Π>��Y�/O�@ӆN
��l
ט2���!��=�Ma|���#��u��t!�1]Y��t����Ϧ^�Q��<�0���xm��ú؈�׻��B��^x��W9sϹ����Yn��["�ϫ��kb�xDx�`3�6��g�E7�Gd��Q�OԼ��l�Ԏ�0S����_ӣ,�ț(��-��8��'?��{R��%�'DA�`���X��*Q��6�=�(�W6�Y��2^92�Θ`/vݍ(m�7O'@���e<�y���1��J�b7l)q���z�vTێ=���]@%�{�-`�<Yޮ�����[-dZ�G`�C' ���^)-(=�dF�h�kȖj��������[J_ h8&��@?�¼h
#�q]Y�6{<4���T�[����\���<\Xh� H�k���!5D)����᭗M�wչ�B2!*
h#0�G���S]l������&���b���n�������k����؛]��2������)��2a\��8�j��n��B�����G6���f��ɂ��ԏ ����J'�me���Qu��)]�|*�����Ae�yÏ�VSj ����L�%:��	я{-�j-��*�@����_O�r�G\��k����pĩ��l��I
(<���2Si�
w�<�Z�bҜ+��O�8�[8R޶CfȚ6ZH�>T���x�!�,� O:u���N��D�bp<0P$���FWui���)��ڒ&�a�U�D��h�����X����q!R��[wy���"��9<6��W�j�sts��u�|���s/�LV74I�4�vP=<�ş���i4��R�w���|���1��E���5�o�`��������җ���准��(v\߁G�TΊ�"Y��oƕ�Cp.̻��{��Q;���P�ы]2��R��gNq:�Kl���@u(�!��Ŵ\/�?;>g�w�NRX����ܲ*���q}�
�8�`���[-�j�2�D� X��;��yz��,\�����������ד��'���W�N���	G�}�0�����=���}H�y�g\��n�p�}q��1/���o���̌�x�T�d��u`&�[���9��s�#�������I}$�RW���Y�qPD��x�"+
���:�J�Wp� ��Tl%]�^�X�Q(�	dh�9�A.�vL��lηjC�q)6�R'��cceB
��/�cц%-�<�oC.O�;�O�M�2��q��^�~:���wa\d�O���E4��
z�B�j<����ș�d���5�)��2b��)K���l!�������*@/���TH��y�%R��;i��o(�>W�<�	���JZ�м*F�P���lm�}H�F����gll��`����aU	�i������>��L���?DwbPN���V�a��������W��`9�T�@��Ώ�B*UƑt,'v��O��. ��k����RX&VDkF��1�Ā"���r���JQ��$�2(ǲ`��:.�'o�����mR`�\g(K^w}]xRN�ZUڻ�˟>�!gO�8��E��/�ۜ������o�{�y��!�1YN�)P�*?YYd<��j�Γ�)��Dx)<)�hc7R@��a�?'��!��	�UA��p��;�B���~��.Dڗ�\��s����wP�����c���FX��~Z7m�a����D��՚&r�,>��Y���'�Ϙ:���)�{���0�]^���# "�қU���Uq�ά�}���E�(:��܅7P"���_�����-�єe��U��Fz+Ly��^�O_�����$P�Y J̲K�9+��TkoA��Q2�U�|�nUb�������ۜbY%�:l��R�?1�����?��}�V�����t2�I~�t�R���u����f�ĺF�6e�q���߈��X=��hY����%����n-h�<0Z�@t��&��?�U�
��"��+�"��{��(��jK� �ex�X�{͚"���Ɯ�ۅ�(��N�oCxK�z�^׆ɠ% �;�9���Ѹ��^2K'5�W}�=� ����;�ݐ��w�T�s�/�Y���}�4��P�dT��Oq���F�]-2Cx���t�XI���M�3KH-�핚T���=�e"�*��M�v�
#��"��β/��k���t*_5�=�:Z�Hb���" �LS���ٲۈ�*m2wv=�*+�, �k�W�r�J}S��lO��x#Sd�ԟ�xY�MwxI��ڑ>�7LHȨ�Vb��"��6A���6Ŵ����w��s�Y����`�`����JP?��U��C,̧pk�9B ���~E���^��)d|��?��B?����-N����Z�L��ڀتP�L�Jk���*��	0�@f�����?,�����))9���8����F��C����^�B��T���ڷ����40\u��-��pZaB�BW�B
&���4Z������%��I����9?%^�T#jZrT׮�8��IX���v�WH,p���j�xfw"8⎎�̙�1�)a��_�]t�����&�s���+\�؍��#�rBb!��v��RJz��Eݑl���J�~�h�;��U�}<�1�N?��{Giӭ�7h��*��4�n,�5�<��OP�P��L�7�8����gs~ly�O6��ym�F�Ɲ[s^N�gH�4̘�~m�Q9�3�o*�0�V7TΒ:� E���Tu qT���j}g:nd�W2m-�cR���%�:����q�V�!�Ib@q�&$�{qC5aܑ�J�[(11Ԉ
�Ԯ��X�n���� �g a!�X�\������g�
Ƕ37j�|2�:�)���d��JO+4�h��R��$�{����}��"Ӗ���=@ԥBT ��GR���$�:TJ��9��@3�"H뜤��h�ted���2ǽQd��K&������o>/����E>>�j!��^k��}�0�Yq�[]���"ޞ��V�C������8���'�gu���H����3�g/
ET��R,O3n	��=�6�8&�f��u%�{��� n���6s]�^����M�������.��@:DIs���S���\�B�Jô�|��栔���|�+�`deP*%U�O+��m�ĥ�7�������'�CY���m&����Zm35���\V�+�I;&g��/x�=R�^������5t��������! �h@���[������@�kr��Ƴ�W�]yZ�XG�Lm�Z�!"���(?#6y^"3$�2�>��)�˽;���B�=u�$9�u�͑����O����_u��C*:s;��yPI�S5��zo�vI�+s��7]�Wk�^�j�