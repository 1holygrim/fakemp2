XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����;^��zm"D���=/5���YՌIЙZ
��&�h!%��'�+���yAN���k>,�%��э-/w=p�o:��XM}�27;���8r�	�U �����}�U�ͪi�L̀N��w�	7&����uaD��n�����Č���B���N��Pj�W�4�X�mk�K�6�o�|0�})嚴PL�~���&$�o�xʂV�#����T���f�� {ﺀ�Xr*S)'�sJ�<\��P��#�`���
s�~h�C]�8�;
���M���4cC+-���<�_��W����S�ZrC�"�4�p*<��Y�r�a�֔�T�˦��vئ��8q�;��x/�-m��MxRܟ��ˀ��~��)ґpz*�X���o �s�ˀ/����u W�A�?ڳ��N�� ��26����@ǲ6�~%�Q}�}��x4N]Z4�,�R;V\��QCv���sbqf&
���= @]�i����A	�U7��]*V2�0HW,F�gD� �ěa�vzI����^ѓD	��f�wW��K�ݫ�xS�o�#gl�\>Mf�Y �L�8�3�9��أP���k
���� ԇ�>q� �0��T�IUM��
��Q�sl��E3�<�*��ŝO}|�BͯӲUB����X1.���rX�&�f��49�b��D�:���e2�ϲ���.��|�
{��GI��JQ���� ��׮���� ���w��:�r�9�z��3�� �|��I�Ϯ���xI�|�%�"��G��@���}�XlxVHYEB    6315    1790�(9�\"w@�����l��IiJ����߁ں>0ዙ����6mC���)T)NlDtR�/��7�ڒ4���"PKd-�g�Q,��~�W��ʚ�*/��	T�-���L4�t ڠ�����ާ�!�	��[?4z�b0�t��[����)0;X���q��vW�l���� ���Z���ؚE��k��Ʉ�T�r}��'�[�5��3�4�fa�E:޲�xB���E�ǭ��]��^"���E6N8��.@��i�u���|��>mN�#�~�t �f��	M+k@[�I�ͤ�� ����?�)sS}9EC��&��<?k���0��y{I���LK��n)۸9z�ݦ��w4Z0�X��:��,[�s���R.�!��m�����������Q�ܘtBW*�TO&�Հ��/eo䚬���;�ZL�I��8��3�NG����M����j��7N�pY@>��H�W����8u���X����o��vAuL��8^[\8�����Ώ�q�s/|:@�_L:�g��LP��K�-�N�/�&��[$��d�9��у�N��e4�|��b�2g� 5p�(@䱴B�	�� Җ��/��x��¸ھ}��;M�2�'�A�uCۧ�l�ʌ�/�SAO�u���Jy9�~�_��
�����!��M�3E&�Osr���q� &ZOё�|H���a���<_��$".SՁe�.)*�GibX�S�:E��8K��?h�������x�@�)*�M���ף`�/�ר9��.���XX:���=X"�t6��/���2�l��A[�φq��Pp��%���XKk��IV����~aˠ_L���X��澲O��}���̈́�rQ5�l���¯�x+)����
��zN�NjuQu�	�� �0����a��Q(�n�^��XC;X�q��u{�������#�?eU]��C�[x�VunE���T=��pZ*�g��O5YH�hF�!s��Ѝ3�V�}�H�ӯ��Y�3���<��ߛ��1�P\�v����Dط�(����F�{Y6��w22�U'W��)�n����e��G-�A�p�#��*�b�o��wZt�o��p���v�*�,�m�Q�oz�k�#��#��0�w��gT�͎�U8�U2^�~����g�Ȃ�e><g�šB�q~�8���&�\�����$f=�H����pp���=��22��L�:�h'ݕ�B�`Lj��k<���A^��������/Ҕ ����2��IC�KX��ɔd�u>	K��-��tK�&������#�(R9�t�0���|��U):�b���͝f�D#�W��Q$Jy�5��&g8�'�����5��h�NT��}o:�� ��!��%�4w
�y!I�R���v�@����: a%�]+�ԙ
��o��B`p�0Zpn[�n�tŅ-s�|��}����ht�(;Pt��o�n�}�Λ[@]�?� �o)�
�l�n��A��w��Uh'���{�[x���!��5�[V ���[�Ѷ���:���,Ex�<��97��O�i��n�i��C��H��#�:!����۰"��,	)g����H!�ӭf0o�X�c�sW�n��y�6 �4\� ;�ZYT��Dp���ۆsՏv=|G@�E����cE�k����o+�	Q��WIE/����(��7����@t��>i<��p��<`��h���Uu:T`�ꏆF�)(*o�]d�λ���#9������Xn���^��uv-�yD�҇�I���([����jH����y�n>��������؉�|�3�Rʾg��ܘ����
���������'�m�.ڰ���q3 �`j��_tǏ���J8����k��G���������R
�k3Y��5�.�9/��	+��3�`Ck�
'<-�;4nEu��ʛ2�wi����>;DQ���)�U�a{\g�hP���-��/����1�X>)�u9�*%�X�+�d5�4�&,�&yL���Mx�h�I�,��G��s��UQ��=����ݤ2q{���WSB��w�B�j߸��`�Q��w�ͯ�x$.�\�P p�;j�>g�~�Yz���~t'�D�i,��T0\�)P�# ��p�ko� ��S�(����R��gL�i��&��,P^"^�viy/I��
&	4�;3�m ^H���4�Y4*}��S�J�M��$l�2Թ����S��\%Ə�mPEc̱p~�����6�����Sxe,�������T���G�	�>ΎTn"�㹲�L��Mp�wy�Q�3\��]L�B�ٞ'�A"�W�O�E���9� C�v�?�}�^���&�i�(e�@����hT��C������\��2뫝f��xeM$� ����[����!�|g1tH4V/2
 �4I�����[k$�8izE?.J9@��ˇ8v�PP��"�[��տ_���B�_h�ƉW�A��'+�u1�Z�|h�ln<jq�ZKy�bU�U�#�������C�(vq&��}�����۸��A�t���#y�����+�{�}ډ��e]��[��D�ԛ�H@a�jw�|(#������t#j;���pF,]��ZU#��%�vsi����)�V.m���K�莅��4*Y��(Q�
�yH�j��j��Ss�k����x�Z��R���t�/��������-�4G���ʝ魃��݄�P���#�U�nW�ٚE�7څ�fuk�V���D*�d�:�j�GhѣWx��tf���;@j�NW��Q��5�uWs�� T������;�}��:K�o�ք�x���&-B�_���К���f�����Ϻ�d`��:/v:nBF��	]��
�-�|*��^�2ݕW�T��XC0Tr��c\�S��8���h����*ڙ�YRй�������O!�z�"�����G��� ��9��b
�,;���9�/qt,�z�0F(a��U�n�F�h���"��F���!<���̚����P������s+M��C̈\��Ϙ�\l) �Z��( $X'WjUbn����B�9�fo���=�Zۄ����KV��L�M	y|��7��V�L4`��c}%6q�?;�p����D�b7�"}�gԟ�]��[� ae'ܙF��2jbؽ�5e�v�Q���]y��7=��U���SJ��x�QR�� �|�ZN��k��j�Eϓ@�w޶�)$���e0�'�2����<�����Q6��E/�w�j�����S����F�w�c�`K|9o&�o�=k\p3~G�(S�"�N[��g�O��O�E��{�טo��e#��[��潷���o+� t��B&	�ڷr�Z6�o̶�}�'<��8�X-G$V+,�a������u��Z�_�?�s�61��<�9%���/(�O]�z��¼w} .��r���p�����w��J疵v� H�_���+�n�?�4�7��!���uq�d(�,%m!�)2.�J�"���]��hXs��b>�{;@��	r%��.�}ҦpJ��6衻Y �&�x��_9r����^݋�?����Z��ɛ�)�Eȃ�o�$X�/C��.����bS�Rs�WV�mM��%�nLi&����q^���1�:�����~w��@�'ٛ=̟���Q���N����HS.�V��=��� -�_՘\��@��n���Z������\��#��f|��H�x�l_ �W������#*�7��QQ'�8���4,l��OZ)��[���u��An��_lG�̤c�0e������,�\�䊲�2ACX�&F>0�Z_N�#�kW�Z�����,�'�M��WۧW�p� �fz��i�}�v��d��G6\u�R܌J���VH�Պe]p�p�O�,M��P�ϡj����n�qQ��]1X;����؅Ag1C&�yqOS�D�g�jX���t�/��ؑB��\֖�X�hi�,I�,Үi�(�ĩZ�[(_����9 �Gz�v�P�Z��1*cܺ�y�ښB���N6������cr`e����ew���U7^�� �&��6�-�I阱L����,��ZXQ��^ɣ��{��	�ް�,����uɵ.��HIčq�6C���ˬ��N�\�ɣ,(f�F̩��q�%CP�v���E�`.�NV�� �p�G!�h �^�_�{KH��^�Sʇf����,��@�	���0�H0��H}PE�����2
��8B2F!�8�x w�4D�z�h%j�8�M��}���0G7\Q���8��xc�an�k.��E0��5�~���I�=8�`��mB:ܞƖc�%lˠ2}����4%!�/�
d�(ˍ*����seX��}��'x;�͎���Bf����:�)�+�P6ܐ�'$p��%�9h���Bق�6����"�U�lz�������񍟦"�pn�#F>d�uN:_�I+��N�\R��ޓ1�0
#j�L�_���GS[zȕA_9�QP�cW#���p����臜L�h!�����T������n2a��?���fxѭFqrXL��	�i"�L:�t�xM�.�P=�����*�i)��)v��-�Ӳ�3�*1�E̥�|���hո�hB�)pA�Rr|�2��^ ���E8�/s�I�W�֫�?T��B9��ǔ��U,���J�;&�����h+�j&W�:��Mk����$H��8=�_�(w��?&�S~NbKj�Vi氏��+����	7 IH�R>�wƲ���:��i�;f�t���!����&��B����G><v� ��װ����G�hML��9��bgR��.�&-gR��v�&W�A��
59zD8�f\ߏF�H�dJR����ڒ���4D��,jz�C �~��Z�9<���VyW�G��5E�Z u5@t߳��-Y�\�ŒiH5'�'~MI��B��C�P���1�BpU}�r��\�����=Æ�kLƶ�%����n2FH��͙�p+\6mm��nI��|
VM�m5ezG.	D>��
�����Y��
|�/ı��^�H�1j���L[�V<�`R1��^8�ӷ��0�\��.D�~������&����cK�@�J��U�K�[!¾���6��43O�f���5�-���t-�Y:k�7�K�������s͉ҩ�3<-T-d����~���r��L�L|�n!p�!�͠�W�@ �D��P�7�躱OP��CY�]�^ڮ�5�1x M�CaQ���|r,��#e�N#�Ϲ
7�Ge(�"^��V |ͮ0�S���x��]���tuZ�rf?_���z �(a�5��1�H����Q���&>+[����qz�H����̘�t��t-�l`)iԥ�DBH��Kv ZGC@��N����5˴R{�8y��>s�-TŐ@���8���(��:������'o��x#K+_L2&6��x�@�;'�+ȑ`}>�~ł�6��>J������I��Uewҭ�-	�~;0/G��ewmu]}0p�:�`�'�Z n��0�9�����v�j�z��-������d��fWQ|�q�F��.�DȐ�ӑ����0�]%�37w,bq�N&>�@���4�I�{�`֍��Q�����RY\Ag��f�R��q{�b���<�`K�o�"�>�͠��vJf��a�w�s�x�>a�x��������e0�j[2K��10ܐ�w6�G ��\���a;����T��Z�۽�
�*�#���/0M	�Q̨"ċ��0�������L�NE�Jm *P�d?���~�c�
�˟=
�����f$��{�iSt���_��*����1�Q�<"�ld�n���.�^��@G���������eݨ��i��j���2 ���Y�d�>J%r`��Ƕ�C{ 4��8.2!i !P��-9�\?�둩�Gme�T��,oi�.