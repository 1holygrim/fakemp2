XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���������P�3\�'z0�����"� ل�|A����V�n�4����H�^�UT���pN���L�e�&�@fZ.�(��.�9(|���HZB��=����r�HgC���
����+>�+�/$A�uu��C��������}��nR؍Ț�y�hy��WZ��n�n'���z���x`��L��wy�@��A��xP���YN&]vLsZpJ`d�uK�	M{���5���������JJ����^"��AYԨ�݆��>�y�[wEˤh�u|L�+g �I������w��ėdR�c�l?�z�D�8�����,�T���9b���#y%m�|2M�{�:˓�/�O<_�j���QmX>�녚G�>���Z�A� ���G��9�t��	�'����?�����$�s�K0,4K]�j�0h^����o�C�z(2�s&M�dS��a3�F���Q{oI�3X4�:�\�ǘ>�[Qɒ�L����*��ۑ�^K��~�0R���YR��^M|B�*�[��h�m�$�*�l�������M���e��Y�Fw��9.�	�����J��c�VwM#����z�欺5��h�*NX�' ����)Rr�5�g��(~'�iG=��I�g���J{��U[�^�d��K���DsD�H=�٘=6�����X���hyHo���M�~��&`�xs���z�S�Z �/3J&e+���TɄiI�i4`�c��|
�5�Յ?+�`���5ә�1��E骙��XlxVHYEB    fa00    2040^D�yd�Fb��G�ۓ�O����/pv��EYoﻟ06"��"����
ף�xnWJ�\\���C��t_��7tB���[r���>���I�Ӻ9����a˂�g�0�5�f��_�L�1m��_�
_���+}&�/lJ�[ټc?�)ˎ�G]<$��Y��v፸�K��)EO������ԛָ]��U���S��tb�Y�Q$|�,#v�ڊ�]"Їt,FR����\�y,
���X}��'4���l��?�.�+��;}�Kc�2.�ёut/9Ე+����p��g��PmYI�9���Z�ۨ��߸���!�\�M��r�z�Dw�]�Xߩ��QYV)κ]�õ� �T��~��IU �)<^��i3��I�3�xg����G|���a;�D�,�������(!A2rUC��_�����@S�?d����v�y������P� l(��o�|���Z�z:�o3=�}�#kEyiN)
��VHS�$FJ�� sH�SZ�1(K+Yw�%��0�2Aø,܉�~�ی��^�U>�}k|x��`q�DX�>8�p��%,����?�X��
�3:�_�Yb�,����5�vBg�SdE���Jft7\��kE$�D�Y����|�J�����޽���@9gՍ
�t/����#C���xnºMCm�o��ȵ<���C�p�{��06&N�6�g�����܏\������9}��"O?47��
X��VU��*lD �X��r�u�4@~����ֆer71쇺���*�$�^=AS��^G��^ �8��H��pFE�C8O7a��P�bD�c��M3��7w��-O���e�P�X��d�P�]uЧ	j�5y##�b+vy��Nm�S�>��_�l��$hla��� �d���J�����M����pTj� ïMr�����/�i����v��6#�j�e�Ƈ��i��m(k��ϩ�c�[�K��B)[	�q�i���
�̓?�|?닷Z�dm�l���aڑ-��p��k�'V75�a�b9��ɖ�q�,J����El�PZ�4�4w儖7��8��ʚu�1뚾:�6�[�ڗd�)�1C��]
HB����Jۇ���#�^F+eդ�Lt7_z3���Σwذ/D��"����ۍ#�}l���%H������j�� /1��k�1R7�d��i)�l�� ߣ��0�E��jl{��kQf	
�����.i��hhQ���cJ[d'�?V�� id]jv�4j|�ѠWu���ӟ��f��Hqbd�43I��S�A���Z�ߏkGd�o4��C�g�BQ�{����;�z@7�j���i'3��E���'�;�wu�6M�������,��X�q�/��E��+5�CFL���D��i����Sdt�E�v�Ҫ��M	���Ж���.��uv����!{�o�C	$�]
����ܼ?:�|N��U�Eq����㏇��ώ�����,T�P�[و<�mFDD��#�R:����b&H�N;XS�V����-�������$'_p}q�2�m���މWQ�Q��A���4hpT&��_j��ՖgUd��W���H�r�0�.oK��Z����e�'��V%��� ��� ȇ�De��ׇ\�j�UĔR�P	�>�t-�hˍS�G����@:��{��| vj"���1.�M�M�OV��]����e�5<Gḑ�-::D����߲�0X�� �:ɔh�,e��٦��Ee�0�a�i��"QrҘ�Ա �2mpE�Nv�|a'�I��L��0�Rv*
c��s�<��Eb|���	n(�O�v�����Xܧ���KSB��6�q����Ia��ꚑ�9��}�v�lL�� �9�%�U�[�%�>ڗ=q��9��L&�EڬDohx�C��t=ؐ��C.���Xz6����`�S뎂�Kb�@��k�tg�GF�u!s!*���1P<E�p~A������Zy,r/=�	��Ƽ�}��4��'�f��Q0Z+k��ׁ b��f���R��
���w��[�Y����#��i�U_X!�%��jN����� ���Qi�<�T� �/z)�@al1�%�Ms��w~��$�	L�Z��侂YL+�]��g	��l�?z��*l�M��������s����5ĉhP��֪���N T<>�Xq�FV��V��?{g�s����g�9J�0r�n�d8�-���Ds�q�w-�X\�U
FL�y�a.�z;�9�!4��$.xR�T��ͼ�Grng-�Q�6	`���E?�|����R����������H�'�S/I��24Z��tW��ej9��ю��Out^�̕���u�☲�,�)6��y �L�C���p[��>S�ౕʲL��p`;<~D���U�}��v:���'I�}�����̬��wk[���x+z���࿀>�x�����L�q`���-�BM�� D"EVIo�ݤ���Bժ�oP�L��Q����!��ĭ�:�ۛڶ1��R��o/w�q���D��a��"���Hؽv���JGú�v��zʴ����/�3ҿ�:��?���ő�
sNۡ��7Lɣ��<�:>� _wg�I�g%W�p���������(ݤJ��jN����'l��j��'��A��]�qv����"�a���ߡ�{«�F�7i`u�,.�\v��<m>����F��?�����뽁ÙҸ�o�q�.�䴓:&�5�3S��zm������d�k��ȑ�e�W7�y�^ˈiE��t���Y�X�~�޶��2BC `��>O�����F^ S擆��&&�+O4Eh�}� ��.{�N 3pH�h���(bu�����]�{O{�xlj�hI����w"<y�9�Z����f�{] ٌBo4�Q�P��ʛ������U��� ��c_��IM�:�=bA����m0���\c�B`�#-i��y�j /{����m��n��;��w'�DJ�nfq���r�;V�\$��1�#�u�~���~��.N
��:� �����4=�d]}���>UtQ���*�����d���S��l8W�k�� U��I�&>��R�?�\{��c[ǎ�ƈc.�i{�v֕��=��ŐwɃ�A��K���B��q>�a�	H��\8��h��BF�r��0.b����1e����L>g�% � �hyF:����$�sQ���8��Ul�t�*A$�A>8?����sa��Vނ��n�'/�3c�h&�z�9|��A!����뺟�1�d����$nY*^F]�C�u8޺p"_���B�r���Յi̡;�GG&���઀qG�qdb��N���8ƙ�̴ht���C. b���֞7�5���0��6�FXj�!�cN����&p1ۻ~+��a�@e����v�c9ҬlUH��h�ʱ'��e^6��%nFq��1,��P�xƝg��0�h�ǒ�@Y�[}\ ��u��kO�5�Y���j�$�P���%K"���H�c��!G9Wq�|EV�n���2�V!W5y�R�Gd���^�4���q�y���/��.2�M!� e���_�#�Ψ9�8�NU�$O���E��r�v�ѐ���hg���&��1$�j|�kA��Z��P���+L5#�#�J�^��n�~C^��Qe�/`�8eX�r���+�bݼG�I��k�ޗ�zFiU��Y+���AV����[��0���ڸ=i&�<�8*�i���g���K���.��e�K="1|4����1@(�K>W�|��ڛ�����%H'��t�6��r�aF���Ʊ%����et�,��So*BM6N %��L�ӷSw5�%ڒ�l���L
�L�mӯ8���Mm�lt���8r&��'���o�L~���*��ؕ[��6~�Qs���	��;b�x�
�T�Zmm�4jб� �v�g�γ��j7��t-�bAj^��J7�	}C%�����k-�Iq�����B�n��P��]�{db���D�I�u$�np#�9@]:&�aˠ>x1��Lwga��F:��B��T�"�I�a8������ֶ�x��.�����hM��}�@�Pm)���S�X�tm�{�r�A���!�I�¶���ĈԮ��.Q�?�"��)y��P�7������WK�x����8���⋤P����h�z��V�3�H���\Z�\O�3��b�[4�i��4b�B��g@J�Sh�]��!=(7`�_C�k:�*���� ��q]ߧ
��F>CW�'�U��~��_-	p�ea�A9�:�����\�jn��3�Z��k=��C4/����}��|H ���'��l4˿.�Y�[�|���/�I�*��Vs`�9�VY|M�Yy���tYY�-RlvT������`���谱�G��+���%�6�� V�!�hFH斂�-�~�q����^Mp�����ИX}5�_�i˩i��x�Q���o
`�X��� �{h!�)�)��:�8T*�8ح:�R�#S��~�"�SV�>*��l��cz�a\H���=����f��3�������P�4����[H���;0�NYΘ M���^�+����[<�sߥ������_������}��̱Q[�mx+�bɀ
�x�ܷ\V�[���	�3*����}���Cܗe7�����\�5L�WG�	�3�*S%A�b�����Hu�.���@��YЫ:OU�8�%�d)}����(�~�*� ��hjnn��5��i��ؘ���M-| ��5�ى��hd���6��>�{UA���%!:�7�N�I.����;-�w6���o8��J�V˙�s��˺��c6�����"�� ��:��_��y�TW/��֪+�GwAf1��! �A��U/�:ܦئ5��J1'�%�G���hb�ϊ�&�6޺m�%\J�	�:(�&l`��D�)����E����C�Y���9 m_�8���d_�������|~������� Lrǋ�L��`�Z��f�����UsǞىKi#/���lR�-��m��~�/d�X�[�
6ve ���j)J�d������s�' �1Ϯe��R�Q̫6��9�U�
�!x���ړ�Z�4��S��B���n��m��|2~_��5[�����&�A��N�H��ǣԏ�Ozd��^8�p�,L��A.٣��MߐvL���lH�>�k�4��&��C�FM�c�E"h,�|��E�(ﶂv����vF�����8�_���l��,<s �\�V��	S����w�U������ӻd��
a[,D�I��OmΫA?tHNN�=����������W��i�e}��s8w�?��$�6�W0�z����N����拔G� P`�H�V�F�́��� ���1�Y�U�1d�����d??�\�ITc�|H�~i��Y�EЍ��JOX��w�t��fh���ҋ��O�a�|3�����h+���7�e�����#w�)Zz����'�'���˂4ƛ�,�|!x���¹������>h�<�����3�,%��X�J7)��Nu�ӵe��҆��wԢ�W�������xK2;I�9g��T���MFbHy��� [6G� 1|�$�&��hd}�=\�5<Q��*f����-)Ό3�RI�(����d��Y�a�'-ՙ5� ,�9r���"��&x�p�BA�Q7ڗH��C���<0��ݝ���d���6��U�9m�>�u�aY���F�*P��.������-�A��=���� u�&���?�rvˀ�:ڨ�0V�*�.�Ǭ�R�y�O�*ٽ�� ���<���W��ُH��{)��L;���p�=f�Ad1�͂�y�9h*�l��I�"�-uI��!�
NP���В3e�_M���n���y���q%�6n:��)��{�K��k�����M�jJL���cn�A�!X!�Ͷn�G'���X8Fߛ�����X�;�P��$���k˙�"�e���#E_PO��w�cg��L#Ee�
w��`Yp��Ezk�R~@��N`�:0�G���jIB+j�StavX;w.��>m�Z��f�I���K�E^��,��~7�/�p_[v���j��6��/��0� ��T��NkM���O*���v،o���l2z�|
L�.(s�z<��TWR@�a߀2���$]��fk@.�_��.����D���ijD���E�m��#u7A��Ԇ#Z���(��x�ȳ���&�����+Y���X���1̈��d���Ri�*��Ų�X�oV�9sȩ���������e�����?�t%�*ȍAlz�Z�)v�1����t�r�-��R�$�-Ӌ�����9�������e�/�
HͶf�IWb:����L:�b��u���ؽN҉*�&$�D��{����8C6Ǖ�q�.<C�A�V`w�#�[��Α����R�y�٤��U��?	�l��W��M�!��_Qc#U1�a��8�LI\�L=b.i���>:��̩v
ޗ
��:����k�5շ�/m�a�w��_!����6f^x5b~�$�}�=ح.C�L'�>kw@�q��ч]t����i&�m�րD�tZ���K1P��`�E»]�����z���տo�!,|�D��nݳtW'¹:�X1J"g k�6%h:�)��8�h/uz�E��UoNv�Ǐ{/]��Q���U���=.cf��d a�ՅaĹ�:d���Wu#���0�q*�;n�l[��x-��2��OgK��q��a�d	ye,���:��X�h��zGo���i
3���oSW�\�����K`�5������Ep���S�S��r�`^=�)���}�*9%�ő��I�:Q��R4ئ?3���l�x�m��sEn�R��37Ǧ��=ѧ�TYd�]�-��wV+�#n�li��
c�w��`[52�_uF�I3-M��Y�:=��c��"`����n���E3&X�v��1*ZC�zyq�rY����uZo���M���Tk#��%������Z�y
v]��&��A��jj�壳~v}2 +c��d��#�|���D������<��j(w,����"���>�kh\U��L�{�&�8Hn��4{q�M�;�ث!��PYc���}w�6��~D"+����C��V�)�>8`m|?J�2���h�����DR� ��.ߤ���i9���/3bϬ�������������~"����)�1M�x�_��v��ES�n`_QxG�o���,y�⿙&f�H���`\��%/�4R{Rߎ<���c�h��2�!>;�����N���J.?|o��0K
�Z�7�KRw2[Ջ��q0��� g�t��N���568�gW�2�C��6ҩ&UiTa�J3Q�X��㙆�'i$2���Ŭo����uą	`��#2$C,.�Zo�V�P�%��6,E3/�����A�j�;�%�
S6�.�>
*�Z��R�|����`*�fX3�U�b�Vc`q}g4A�t��_�ކ����� r���N��@w�y�h[�t�C�}U�0���k��0�.>�����
�0�Wr��������l�7#�=D{-_!��O������	ÙM0zV�V1
����͹bO��Oݤ��sf���w�Mu��D�~�J�f��T#,��&O�`��9�nH��o�����+�*l�;�h/���Lʥ��_39$�^b�/5/�!;x�1By�mӆ�[]�/����y��kk��Ϝ�/��d�Ą��m������{��DN&Oя�A3�v@��ې"�%� U��PTz0�k��a[���A`PrCI��H�ZԾBn_6��W3Þ��i��W����!/b^�[v�'[��Me�ND�S.���$�c�P:t�4�8?bW3|����v���b,�����i�ǳ :>���%A�*(G`n�_�}G�L;(N*�@�[���3B\?c6y�@�Fld���4t�6�ڃ�WKN�D�t'�d�ܐL���t���V6f]�8��ԇ`g��r�%x�-��*�Ѕ���#	X41��O�:�%�g vK��I�R����߽,��[P���'��\)������&���;2T�Y/�M������r3P0Lz҈#�K���XlxVHYEB    4f62     b50<�q i�"���Y��V�B.�Yr��G�8hf���_8.y�~��(Tn��szH|�oe�1���!��i�v<I�j�V�eo��U�ʔ��0[�'��Э��췏K���;�Qkm��rj`��d�8;g�w%��4��M���E+7���>�M�N#��-�������MR��M.D������#eM�8s)��@��Vy^��L�%Ď�
M��~&xe�&_���&�����V�H�����B�V �*-�����S�(�+��>�S�f�JG�+�����9d�6��(W45^��Ώ3�f%�g���/uъ=}�IM�+����䂾����+L��PK%�N�W=����]�^�{����V�w��d@�:cF2��3b&*쐄��U�ަ!Ȇ�⿛�3��Uɨj^Ƅ>x�n?���16��N���F���H��u���P�B9d��z�({=
@�7F�{�8v�p�PH��G����r����9��]u$�d���I��NE�T.j-�#�����&��\�ͣr�$���۳%���;����9��x���j�3�d35xw2`2!0w�@Y��=��+o�:��t�w�P[������C����X�xv�:�����L2b��w��o-7�ùv%�'�=�Q-�\V�eN�s���0���! h��f��l�J�۰H�p�ޝ���Թhߒ��}p��&~b�C'%7%��x2M�T&�XY�c��$�GR�A�x�~W��2Y8a��#��.�0����p�s��q�Q���ۥ��p0�w���wcT8��"V�t�U�q�W�w�e=�"˂��
�.����@��%����
��q�	������o��O�C�}�� �RK����]�	̱�D�?�3��M@�����o�#[B	�d�۽��Y����a�i8�%�<m0��6��}��f�};��S����kw
.:��y(%��ljR�&f�S��-֧����[,D�F��Z�S�$���%�/3�n�iS��F�X&�F��2�)�t��'�K�ɩ��'A�pO?���L���r33�A�n���:B��̈́���*�&0�L���!���	ڊ�h�E¦f���M*� ��f�J��#�|^�~Km���#�ߒq��H!�\�v~͝,�9�`ez�a�Q��V���O��%�=�;X���I8�!�����$<�4���h�ceX��߮�H.����"�qRhӕ;7́-�z�'⾽�Np�R� �`��\��1>CYB�9��IK�z>3M��>��q��� ϧ�}h��s�~�@�ow�i�7�f;���g�i5'_ӻ{?gL�����'�m6wL�L_R��V�$|w�5�z@��f��=a�v�Z�\hA-�$���6�.j@�4;��g�A��Q1�y���7{T?B��_O&n��}����I8�w[�wJ��[:\&?}����ݦ"D ���Ȣ�;������~L!~�`vU��:�K���k����"��$(;}&"T��ĹL������L�s���m��D��
�'}�%/�J_֝��|v�_��Hב�q���(6�}tl�-0��O����@�O��.���q�%�������m�K茑T4�Y���I�1�����}�s7>P���AhG1�<���t>���?��!���W�n.� Pi��E���~�5q3>�n�=��_fji�iu/ֹ����Nk����k��
PPErg""�?�oY��&u�T�_r���t��m�K����w9&��m�j�h����bj��ġ��Q.Ȁ	�uM��B�);<V�'b�Ql�.�B|�L�J(�J��2F��k|�O��@5��*`�^Gs<�x@�-���= 7���96p�Ťi�	0mVA�\M�I9�t�X���5;��m���`��[s𲄅R=��{C��~����LkN��B���º��5�#�P�G�Y� �j��'Nb���=0c�hU�芑M��?ۥL�9�+��fx,��x;�8P��?nԚ��*\)H>)~�q�����p�����ɹxǮ�/�뺿I��;��e�}~=�s�'�
�i��y
�ێ��p��|���{*�Z���^܏��ܿ�a#(�'������?٫ܻ;���tҜ5����Z��U�EP�lܙ7m���׹�c��C���*)f¦�`@��Y��F�	������]�(���o��_(΂��>?�;{��+ڀz1F`��t�o��Owb�!�8QaI�<�G�B9�U���	Va�� 1�e伅%�'��͎�m�S(8������=]�	��6�5CY������sz�C�\�O�J��&u1|gPP���.�Ji���h�ƨ'�v߅jN&�.�ܯ@�t2�M5�3;��֬Dq�u-q_z��f��C[�v����x��r��u ٍ�W��������?2�s�D��n��[�~�}���8���O��W ��CM�`	xt��y�ܼ�˫=�O�,�r�q��b43v8��zQ��4�YlVXП�R�Al�=��H��W�6�RDCǽ�'��l������x~���o��tc�x��?���RX~?B��U�,�P#�S��1XXp�d���E �������SRB����ph��B^���A<A	r���u�v̛���MS�>0�/F�C�͝_�����Sl4��s��(�T�-)�m��/����c!6`K�:�|pA���J�9s�l+�@�ZV;i����F����b�Bc��ݚ#U�I���}G�g��7O���}QqN0��֢��SJw�3("�f�{�6��Z�xL����N�T�6..Ń�����P@�y��K�*�l-������o����6Se�q�