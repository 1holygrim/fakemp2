XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���E�	�����rz� ������(�+F�+��n��pR���j���/������l��t�,d�;j.��Wz��f������6@�-�"�$C��Ź����T� ���*.+�`?���s��p�o��8R��EE�L��G�,@*�(-������9��\փ���1N8GI���-��`9����t�D@2=4������3掀�U���VJ��(����mB'�ve�m�2��L�����y������h<O�Wr�{��ɤ"_9�F=eY�*�A?%<�
���4N�#��K�B_�`x`ܪ���Wh	���pK��M&�lG��o��h�a��8���y�C_�&�1][ȭ��4����HTU�$/��������X�*�O?��17�ffM�2n9�����+�h�(�w�ij+_a@�兙��k	����b�b=���\�@3�\̝�J�?!1ٵJ��X Ԍ��uZ"�ћ5�\zn�T����5	#��YV��V�rǇ3(��J��A�<�
�������1�,�����f�q'+�{�t�,��"��pSH�M���Xiϰ¤�����gI��ߠ�	xc����p)�_P<�O'���&=c/j��g������ɺ��i
�U/BH tɳ7����QF=ѿt��;�u�P��Bf�?�?,>����Re>`��@h����݁��w�?��h��-/��.OM��-�� �@����؂��}���tj'�����>���XlxVHYEB    5fea    1830DK�^��L��p����A=�e��6���=��zЇ��% ��B�w��孊��&m=z�=��,w��s<��� K��	�9�-�mx& D���E5�������XL@q�������/�;3 7���ﺱ�"rDYPa�қ5.��8��| j��̼�oV��7�&ı�V���.��pNl�.��_+ʩ/mZ{�R5p hC9c�i����ߥ��ԫ+p���{�B��آM�|�y�K��ma����*��^/�w1<5/\T���0P���{���+wM9+��r�U�"\2��z7s��lpd�s�S��@*�&.Az)1;Έ�@j��C�M�9U�f��5�Cn���uAI���$+�m�&�@cT��b�󚁎M���O4�`��>��/��2�̨P��f��B3��A��3�=DM��� � �'A�'¼{��rcF�� G.>r8
�8�Kr�c/�e�-���bZ�7k2����y2Rb;`��x��J�M'��_!^s���sRafb�F.�x���;�O��wv�DnW�3/�"�� �Ks6�����
�0�`��%�i}0>�,3L��tJ�hnMth�:f3��`��E}������&��6vi�GY}��?A#S��?ž�v}�g��3���ҝ 4$��p��i�%���~j�N0<���*hū�m����Mjq���EJ���Q�}R!� �b���ݛ�9�>�%����ng�p������>.]�Ѧs�#d���¼W�;j97&�Bnck�۫�*�4
�}��"q�7�����3����lp�xk��e�̟�\h
�#$�fk���ܠ�%�>�b�A?�7�����C��t1a��_ea��lKܬ�a?>��3�YW^ޖ��4����u��f����������7ɽ�%LU�]��Uח�5.(+�%Iސ��B6|M�.����ΦQs����r�͵�#J���d���%�[6f'�(�Y* |!'s�^�%I��C�TO�v�҆�����A�D�
�\�+��p�����z]����z0�b39�n7]��ݴ �zP�g��5 �wGC��\0��]@���Q�rJɯ�c��,D�]�N;�*��h7�"k���~���\\��R�~ ��~�X����@�i=��ԟ�x����,�LbPs&�%��D!�p���(�L7�ڜd�GHbm�N��MԨk�����q9�M��!�^i�!i�y`i�g�w��FQ5dB;2�������v�q�nAZ��b���:9�%�d�����ukld]|n�@!�����F��3����xT���~IXl,��.�`����TK(�=���٠�b�ҡ��gl�DQ��d�qXd�:������nt��V�5��4!���ۉ�D@����z�P�Ù��橆��D2v�)S{�>V��"��� �A��],�(����NReO��1A�2+}�TxP�E���kN��9T~Kn����+��]��&����(����O��H��3���O��ZԜ+��q�������V�B9�m��hz��5
;��w��8d�����Se���"�t�}vP��<���!�=������W+��z������f�qua�(T���\T�<�͗"�V��hP�Z��0j`Lc�:[�p�KprE�Zhj@D�`P���%#9�TN�����0eC�T6�$�̓E_��=v�:adN�pܽ�3�J��2��|�ɢy1�9 ��j!�mFW��"!�y��VBJ�*F\Jx(x����|uC�MüBN2` ]�83�HRΩ	��]%~b���0�RU���h���Mg���T�W�r�?x��^-�ҟ�wq����^�(�qQ� 4�P���	�@�vL��J�G��Ak gYg����3�����G�]���ݙ��Ā�k�w^\U͸R�e�0R�">C�0�v���g��{����L��*pϜR6��MG��Xk�5��x�\��܆��r[���t����X�Z �2� H�c�ȟv�;0I�跶�����>�K���C�^����q֓�g�M�	K�P�:��)�e&]ԅ�w�^Ӊ��� �d.a��E3���o2{��I�Qy�+��,4��@�.���Ǭ�@��2����>C���%ȿ����Ji���_1����v�͆QF�����L�x�����(aNz�j�M�4?=���(�S�S�-C���u��W����N�^�)�U�.(��&�d=RS�����jW��W�.���k<���S=���&D/�|-|�^oc����x$��8P���!d��ʙ�p�z�-{b-�gxg�73a�o�0�gxY�5�j�� WF����+�3I�Fȝi�a*My"m�&9V�9�3r�Ui�뙉],����(���4�G	Y~��,+�Fi�+PT��X5<��6�1��}�����:�J�׭�!c	��M@���F̷���ꁨ�{k'N��-~��'�7i5@Q����`(j���叺YS�(Uv��l�����A޷@ZM�|��C�Щ�jn���;^	��(&�1��������_ͭ�Q�[,n/p���a9�g@gLe�}fo��zG�+������[*k�H�����I:P3�Z���W~z\��\�-���!̬�kփ�~�A�S=�V�,�)Ҫ5�k�@Lsh���W>#��úx�v��}j�ѫ�iJ
\�_�9R(�(���w��Sb�k�2�ܶ�ؚ�g&���@�T� ���*�W�/��/�V:�ٜ'�qj����J�izЍ�gYkt�����f �����"Vm����J��%(�J�AK��T^Z���Sw��gh ��<k�s�\|��*��U�,�4��Oba���n4����@#��p^�`y��y���U�F;Hh�J�G9�<�[~]�댱��3�C���)�=���O���ԣM�����T(��,��U ��m��� 3{�D�(����E�*���"����芊Q�lEta�f+�,�Q~���C��D�:��d>���u*:ё��>[k�������	����N2�T���l>0��ܮM�����6�C77)&LY���A��|�F�N�Ұ>�>U��WT?�Y���"���*@�����S�����B��j�2��8���矰d���u�y�u��W܌���]�e�G{�ؐ�P�ߘ�!O_	yN��o��SY�PʶL=�p>"����V����+��DW��enD���ˢ��5�Cмd���=�7���"j�� ��_#�̈́@Hx�>$%���*�O(ź�	�T��%4�n6��5���W��W |���,W�� ���L�]�*k��n�'̾��	��ʍ`v��|fLG@�}�+�kߍ��>hz�u]܌ؓ�ȘhG��v{�g��XK�՘��G�8{Jh��ƿV�"hƛ6�<����[ZǊ?���Į�2�RϛNNx׶!`0aaV#��m� �X���N��b�yXT���0��Ñ~�5������UoF�˅5��tcZ������h��pK�����J+Q�ـ�h��haޅ�tң���uTds`1�8��B�v%�eh�_�lxg#�tT���)26ٲJd:2N��>��U<^ls���ǑK������G^ꐎbN>�<��%�ڒ@E��.	�1j~���X������^��/h�Ȝr�`�c�T� I�	�il&=���n�BmB�!%�=&��u���#�k˻b�0�i��އ��]zl�@r6x�=i����T�0@�|e��@��!Ø,jU�K�Uf^2B�
v+�-��b��%m;�{R�n�#�;;w���ƫ��t(���e?
H4�L]y�	]���N�_���<�~��u:N�6b� %e�\��Ur#���`�N'�Kh�-��7�E�Wkѵm�_��W{�\���*Ł>��m���싰E����x-{���q����Y��E��q�\��8}"�b g
7�&�����b�<�]�.����a&��ű��G�7u�#. ʟ�e�ώ�z�H��~�0�Bկ;�!�@Y�� �67e�s����?H��YhE6��d��o��j	�T��1hl� F �@�&K��֚j��1j�c�d@��O� �wS@~\��kqhL���'�&E��|��F�J�/*����bҭ� [��%)?��a��w�x��ڋ�������4���4(�O)�2�6� ��P���e��+���H/k�6��gS�h���t�c�����$�c�}Eo�)+�����ƅs޽Zt��(��ʗy��d���d��fҴ�kl:���6�U�*��E7-�E���$��p��RM���~b���:� �Q�E����|t'�0^~���gf��2�$�����4����>zd�P�=~�8!��j�
Ԥ��F�����POٺï�W��������M��������l�롎V�=L��SA�Y]Ƥ�1��xύ<�%�'~HZ�"���s�椥YU}�T4����|���\���%��A�l���� �,;�O���������l�����ϒ�Rt��%�#2;[}�_<�IqGU4ߑQ�*҆���/�>�"����@���� W�ߨ��|FLndE�cr�N��(�*� :2�E�H+3�I�m%
�0��/$%�6��u7~P��:E~'����U��İ}�����[��A"�.`�g���-� �g������'�B�"o_�s,n(�ă�S�Zބ
N@�ȕ#�?M�u6�0|]ȥ�C#�����o[�`^�\勘���{��UIKϔ$c�z����s�i���4bi$-�K�_�E���m�<'A�W@�N�	�����o��U�!��mME}�S��v�lͅ�Y���>)��ǜ��Hht�5� :{1*����ۜ�:�]2�˔� [��]�HXQ i�0��%ԍ���#;h�U�M�=P�5[�5*����Q���$!�]f��e$?���X$����:��c�3��wӌ�5��F]�\�/��g�S�%3�Ĥ��Y��v_v��${���9ڛ\���(�����A��u�6$��e���B?�k��D�Ui�����p�sb��zx�=#a�30��U��Û��uBv��@�B�V�ć.b/��}4�lJ9z⼄�q�N~@��m#)�]�r{�����ӊ�0��|�(ⴋ���"�Lb�g��)P�;I�'��t����-fp�"�H1�07��E�M�G��h;ϼ�n�X���~U>P�%��\���!�z���x9/�*�l�B�t���J�~|��K✀�XZ?)\�Oט��Uq
G�ߗ'`����|d*k�k����1l�ꦗZ6ޑ <�k�+��<�`a����n���BZ�yo�tGEk����Ldc��n�H��p(�e�5/l��R���*���W3Ʃʇ�k3��(�nTx��()��0�4�}���t>�EۗU�/�ۑ_dp�@sˬ(i`����2�z�t�%/ۉ�xr۸ĭ-T.�ևO���6?���oaL�p�[������[��+e��X�����.}����ɼ�$��8��gm$�������ʹ����Vʙ���+�Ɔ5�@|mLg$d5�>~9�^g��1��X�V'_u���R%6���/�*sҫ���KZ�R7��򄅗3^�sQcta�Z���g��$�J۶7�P�@4Y�ߙ�%z�w�EIAtnR�~m�u��~	�&��Q#)lT)�?!��i�z>��g^��a�U�a ^[�l,�$j,f�Y�%�p�e=��oj�c�n��8l�P{$����&��L���?1H.E�5Rہ�Ʈ�� ܃��A�`ª$�(W�L�.�<(E�7�"�4��d� �JC=��%Ƥlry!&J�z�!4tE@�՞Y �)� e2�n��?�%L҈��B��U��n���r��x���o��b��������/�H�xHx��,]z8W�׍g��5O��`��6.o�eRt1`����)�o�¹U���:�6`N���@����A�k�"�Ԣ}�H1�C���&�։D;����\�َ.�1��`��