XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���txzx���3�)<
�����^������͎�1]L`�BO�~��Mte��ҋ/�&�22����W(_m��j+C�����$���;�j�2y=�g�`�`}�gh$aJ��N�d�owmN O�1P����!2�ǳ���%gD�{�D�ǟ����6���ue�ݭ"�ZJWI�+^�+!M+�h9U�V��[��D�?w��~�Q�Ѕsj5��: ��T΀����\0�e��� ��^�z�g�T���UK�T�~�u'��^6�!� )��o�E�I�r�X�x(�
c*���#�9�x����q��P�h��Kw�����&�L��©f��q��iT�Ϩ�	��c��ե1��hx]�� O'N��(:t⨀=x��w
2]S�'J��L!���Ho1�7�jm"M�C����"��ӡXO�����+�q[ ��wv�v~M�S2�+E��Ӆ	?'��#��ù��?%�2;�;�F��q¯��1s@ĕ3�?4�(�
vw�z��0Qn��"�ꌼS��c�=6Sa�/�zȮ��0����f�����+z���b:�)v-��h� �����VOpJ�B}����A�U�Ncλ/A�	__2ԐjOf8KM�#�Kr"� �&�Uˢ���`��jK_*���#���G�l$���h+?���5rJÖ��BB�.��YX~I�"���p/v�:!�w��F��6��k�
/	x�������I��P��Vb����;��ny��C�(@E�"o�"�XlxVHYEB    3e93    10b0$� c��Ѽ������$2<c��>�+�e���~oq�"A�վ��羲zN��BP�!K]e��S�+����7�fF
��ȋL���>�1�H���K�{����n�Nt�4u�p��4R^zv�m�(��v����Gm���n�T�i�<���[4*�a��F@�ɮt�m�I�jز���q��n:u��������':�R���]_�՝F2�la�T�q &��XB����K3=٨�t�mJ9��1E�*�����ǒ�L�;�1��~�"Z*e>V�_�w�Fm�p�`!:������L�э�f�J�@Z���yN���,Ti�ɍ��������0U���` �󞐜4O ��E(�e�Ȫ��X�
�U���&�ԽA���J0D��s;����x�W'�y���y�͖T��+��u�,eyj	��N�KA[�Uɉ���h�!ʆ,��)�e�0p|��K+�Z��?�
lJe� d���G�����o�f�r_��Xr���Ǳ������m�Y-5��e��)W���!��_��MN��l��1�X�o<oM�,�ƙ��(�.aB���N?�&
�!Rw���_b�/���ֺ�a�El��!�v�P���t���Ɂ� !4��.%^� k�"8(��������	�o�R�?¹�D�%5�w���VtV��-�aGB���(L �S��T^*i�`�:���WU0X� l�5-��! �{��z��Kv���f��:(4p�79�S>*�P[P@��a��NdAX�)����ыC�&ƾ�P��o�s�L�'�����\T*����\򤓸�x��EG�����۝"�$R�(=p�u6.���,oN��X\���3�b�c�3��&g9TF
���\�A�f���d`�����M<A�rF�ř	GY��I�0��a�O�P�n�,1�.w
3,��o�=��βafV���a�l.�H�.%~��1~wUpc�MAmR �䑫�
�ɂ&Dn&Hۘ�}.�̿R����������<�T�dHz[X�/?Ъ�K8��W�KF �
	���d'd 2�F��Ye������h2׾��x�P|�ă��)���a'�ĭ�BH�}��[�&���k�GNDǜVq\,�'�p}�#��X��3R;�gV� ��S��Wc~;\�;�^�/�r_�	���I��jN�v��ω�q#`d�se�d[���1�c�輸�F���~5�xP̙H���J��1��V�E���G<(	bm)�v�*u�&��_�3�C��;>�,�6[��W�XiQ �"+�ua�3���H� iJL�A3�Q����*;�=��7�܁P_���pm8���t:�������H��P���[�d��N>ߒ9���P����/�X�׺)�0f��������f&�|�*9S�L�8���2��D�Y�1�X��6��w@��A[��/��P/Q4C#��c���9�G� �Uc�����Xw}��ݙ�飅[����߷H��}��b9Mn5}Td�v��M�F ���M$��O���h���{Lk�3j"Y�Yat�Wߣ��r)��p�.Ѥc�e�+^=�io2I�@(CXR�}g��� 9^Vq
M5%�@�H[�U�����d�(����ʺ�4C,�|]��W�œ�w�<T{��k_��PcL�P�[��|	��2�������R�=l/���}vsx��u8F�gqj�tx�9<�3O{���܇�� �s�����c���)׳���%`���5�*:Ko�~�����m��	Z	����/�K����D][L5׭-ټ���C3.�/Q�v�P��\&I�5��Ot����g��-��G�f�"A���SLA�O8\/�Q�������	��EQ���q� �\�NT�;�囔+0�w�T��j��Z�6��/)�R�2��"�I�W�Ħ�ǣ�{�,�Q��v�g�
�� ��ͽ�����W��/�U�S����Ț����Ӄ\ʇe2+���	[�r�	F��� n��hj���O���qŭH*��k�У��~�Ne_-`S�ii����Iu"��~�e�P�@r�g�Dp�����?���}��~���p���B}8-���$!�ސ֑�K���o��Ƭ�,��:)U��dHj9y�pF�O���f�����ϬgM��8p���L���Dۋٍ��	���C���qy��|���)A�}M4�Ġ�8�fZ��6��[�����9��*f̰h�F/M��`u$��Hr5��!�C�H���gŴ9�*�'!�*�9-&������3��g|����? �q�����k>h�/�|Ev�)6�i\��$�lPaQ�ęi���Ej ����䟍������Y<H���6sC���r('� �2�ߡ�ף'ta8|�${��s n�0	�V�)��A֊�{��&�[2�����!op���7��AFLs��Tn
���+�8S��]�{h��\%K�]��WW�]eLO���5_*Z�H-��+<��D�f��z'������{����U���J�34�&�ѕ�����5�p���Ȑ.�*�>E�X�6�H�@��1bP6)�'(�3E���S�c�	��	����u���[��P:�J"�P�k��W��d��JD��-Ն�r�פhߐXJf1��Ѽ����4j�c~���K����gal,�Y&tu�\�u�����#�/�O�3� �NC��?h�;���sDL�}���}"H����NH������J�C�&v=(dߐ�8�x�$a��f�W�A3.(�`�L�~��p�R� TU��G��|�@��m�`]?1�M����UJ6��M�
+5�#ۗ.q�g�n~�QR"��z�w��:T�w�e��+�zJ�H`��q���������T��0^D>bn����r
0mDcV�ɼh��>E���#�b��L�}S��h�i̺��k{y'xE��\���P��x���8� SD�\�pp^*A �~�:y���6����	�Q�|^�4�d�d�v9��jX�@�� #��C�^��ā��d�@k��	9Ι�"�k4�c����=ɤ ���ٴXTˮկ��V�o�D���<����7��}��,��q�[[�7�)we�l�,�b��h0��0��>k�U2���T��?eo��{���{��&�*�S�Y��#H��I%�qU��߫aS���PR�Gv���*��"O�x�s�e��2� �c�H,�,��0ԎF�!?���͓m��l�ʜR0� ~uή�%|R���2}_��OܧG'�H7��,�i�F��*����X�[o��r��VZ ���Ɍ��*���Xu-hW�3lQ�jC]'����t���c�')Њ��+t=F�܃�n$A���HJ�����:9���OibyQe�Z����U`>���S�q���Ζ��b=�}�݊V̳��V�9��ﴧ��	���Ȯ3~����'�U�k� JӐ�eV+�T�mS���d��c:��=H�99�`�/���b��=���TJ�o1?�v��XB�eз�<�\T���M.avdGw�ӳ6{��-lB��`�RS��N�=i���5�����C���?����U3XÃ�y���*�A+���)qL�����5q�_m�9�9�e�:m�Һ�EL}my����Z�c�L�Q�7)�Cc�x<6|�
w4&�s�y�x"�J��>�1�t+�qm�C�@�^�%���EM\Y��9�|��
�F ��R��,5�f��u2fh����:X�^,��p���n�-]b���o�t�қɩk�8��?�>-N�g���h&�;{����S$��f�'A'|]_@!� �G�]R��1�l3�H�/d�*�O��Ew<��`*f�3��w���>��T�KMLc�@Aѡ%IJ<�_����'���g�wO�Ta~�5N��cQ���sǹ�[ߖu-1G�6���^�[��G��'�,��ʿ�^�ɮ*�a9�
��g�aޤ��nY�Y���|�Jb��l-;��O:_[����,����>Texm��-��֙?	r�u��l0����;�8�~��Uf��..ă��R���r���pH�.�V�Y��9ʺ�Ai �N�������v�0
1�Ϡ}eNEf&��_�4�-��=�j%��{���-=fV�h;I�&�GwG����)���r���3�,]&"���
��K��C\��͔��ʧ��肑0�+�)%U�