XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��-�n������2�n�Y������7�88��$�����6d�`p����S�F�<��1\P�^9x��p@�d�uBe��sEn�e.�u-�@:�;�N�2�o]��9=gYF'J U�$	���D���W�������J��׺%O�>IvåyM{⠃8�-1��m���r7�p�cd��j����aD�	�o����9���Բ6ʿ��|c|��E"��g�3�"��p������S��@:Eg�Ԑ���#�6js�u<���gH%��
l��]�@@S��V�S%���wt>�wp$��]��-BX+ Y�=I�l�{׵�����`�.��+�}�?������>��4���,��ꧬ]%d�Ǎ�M�����lɢ����3QA�?a�����>�Ai�*��y�>-��^�����O ��t9ɯ�^��5橽��|ƛ�Q��§�3l���Y$�K2�5�z'-=˾��dkav��t�b���oAc�ԥa��[��\������'Ne��s����d�e�8CJ�d����쁂<�&��x4���1Z�tK�A[/�KbR0�h�u�,�+�I�R������ˍ0s����`O%N��2|��7�;�6;>�jn{FJ��GCy�Z;Y^�/<���8�KA%��-�@���[��4���+X���J ��#&��R���hu����kS}-΄�eʆ��'���g��Pö�R��q���i��z)BB�����X7�ViT =K�������kkc�
����:w=e$����:*i6��
��M�RB�XlxVHYEB    95d3    18d0�.^h�5��h/�yr���_`P��{i���}��ƃ�{����oU^�w�`��nx��vdǕ�R`Qf�Eӡ�1:@692���)&Bb�̣���V	�$;6���P:�I�n��B_I�r�j�_>l��|Dv��:^��Z��$ѢUE�_/_�"S�c({ly8{��G�64��)�K�7bH=n}im�����k�� ^��n��tgF`o�4Q�-��N</�g1��-�7= 8ѝ�Uqx��_r\�V�X6��W��l�m�ar�����Z��y��@pe�c�F�����dc�X�����BDw=��4o$0;�1>k�'����?��p���=��V�5������������
;Q
��a5�0Ƽ�'&j���I.��W5���D�?|;~�V&�]�-	�$�RL>�7�!�@�� �FF�W���:^����9�$��3˖X���0f�)������敳|��m�ꇕ��1#�w����ҺB����x�J0�L�k?�dN��zN��İA��|	l�ň�o��I\&��֬߰��-�����2�&"2ՙ�4��S�fx��%�Cwv*+��8�~�m�d��<�JaR����T�gt���)8t��t�ܛ.���Uz�[�9����ݴ�6���iz������#�ȱF����l�[+\��D����\)�S��bw��G�Q����?o����b�d� �	�Cf��vo'l8����a��>l��/1��t�~E��������j�t�$�&�U�˭S��r�2횛���+R	�n��k��Y�8R k���iqˌ�z(���R��Q/!�����ď�C�y�K)?��w�?e��Ɋ|����P�N����_~������F�~�w���QZ��{�%M�:�K'@��FPr��|�(��ts���\���(��rX��v��;ʡ����Uw�/-���O�'P�?�'6>��kJ=4T��˄G��<�
-P�@��𱙅�ǳE��-���T��.�}q�%B�ݿd�/�������<�����	z�-���F��V�oճ�خ��[�7Bo��D7�m���7�q�.s�8g���}�KBzT�F���H���9Z�����KO�v'���6fj{�|�{����fu�w�[J��M<ROm�1��?����yH%$��_l�����K�xnq1v�b��G��My��j2�x�^��b�& �6�#E�2�3B|��Y�����[������T��S,��s=��C_:k�4TiUYQl�.G��nӼ�p�?�� pʭ:F�_<NA������Ky��F��'1@=g�&�))�$������g�<Z�q�{ƾ/`��!$3|��н2�^��Q���Dn���:�sO"��� H�5"e4fM'�q��B�fvQ�:NP^0��FZ�j�=��̉��N���3�F�RG�	x�c�K���t�f���+����u�4OЊf���u���5�&��I>�Z�뵺�d�0�P�%~cs��)��Y�e<�3q��Y�<0M�
��DY��[XX�,+]�N��1S���+Ґ�W#HU�K�7|���+����C���~)9B���FYr���5m~kF�GI�������x�K��5.�{-P���g);���yAz3�`C���G)f����
�u��2=X�/�o��v�ǐ�#f��jZqۻ���R�x�o|�}e� ��-�T�^X/�%�HU'?�����h�׊^�� �=���V���,j�Aq��4�AT�T���2n�!|�nKG��8n7
e���)��͛ Qp+X��K^t&T�(��e&��*,8	���]jYh~`�ؘl[���҃:0D��Č#�4}����\_%`*D�˽�/���O��k aom��y���Na�4%��]QװL^k������8��9\����ψ�i���Z�(ƫ�����q��JjU^	�L�Hcq7+�����$� թ�V7��>���푓�U|QďC��o�@F`�V�A�����kUFL=3��"46�G@��\�Nt�؜�*���4&M_�<�y��� �v�G2jQ��؛U�����GX����y��r�%A��)U�����^���V� *`d'2�g�%i�a>�O�jKq��ª���c�r��]��]�?H~����T3�V'��_w��4�:e�8w���0�k�Y�����p."���v5�NؔYb�鞢q��tP�2f�S&T��	��n�5;�z ����p@�9Hϩ��� p;�)����^{3��C��������TȰp'��_O�Y-�Q@�����dI?A�� ����#�d��mE�:Ӑ���9A��:V>�{�~�S���o�t�Ř ��!��KS���2�\�!�t��E���G���!�*�߷
����
s+AUh4qR;�� �����+���&{&�f�:�#b@��	~���&�2��lo$�zWR9	�3��ػ�D�#,�"H����R��q[�ɒᥣ��1kK�ng�^��.���@�i�p�w�����F���F}������\����q�o�,Ǔ�w��߸�QH[A��ex�
L�=1��@��MsR�4���n��I��4�����S�jD�ŭ������{��,�$�o��4q�$���8��kz�O_��h~$셱:
��(����h���%w�a�c�*�]xLy,W�EI��0�_�	KH�rK�����t]�L������FQT�좡ς�9eY����,0�1�b��^|��+��W��:�*<9�ӟo�PnJr��O��;�=�~���}g�i�y�B�JR��0#a*��8�L�}�=�pCeA�k�(ho(�OR&
˦����n�T��8��ҁ=уj�n5v��Z��a~�R����y^�<h��:P_:��Qn���,�����+e����m�F);�l���7��M(U���Kp�f	�	��9x��<I�8���䇪�d�E2�Bp(��9�(T�J�iDP�Y.�9��9g)�ry��l�N�n�Hi��Gn�o%ۦ�����_h��bit�H�pŧ�5y�>&8�R����`C��'=ZՉ���?v��~�ti.��վ�ʐY��d�O�O]���X�?�qJS����!���TLOS��6�U�x	� ZDq���ϋ�q��t?s�:������>Up�%�#[Gw1!U��J�J�r�!P�Υ��gy7:<�/��h�?'��m����,�4�O'��9��%X$`�kW��)
�S�50��ɝ�9
�F�j��*9��A/D�/�ow1�ȉB|v>j����.9<��~e5�؂�����C��������\�l٣S������
���5�5q���T�W�.����6�i�y��k��һ�]fw�B�n>�Cve!=;W�x���]�,��َ?xQ��C�������}y�s��l��$6A�[��y�wx�eѯ�$Rr�cT.�תY�l�R��6�g,)Gs�٢첾�mC~d��fQkS�fY3�jd�}{�GN�a��:)D=`:�2�.G�;�ys[����!��HD�}�ٲve�C����vN��c�~��Y�ǹ�G
#�Ł�<�'ñ������sy��߅,^)PR�{�7���`hEa�E�B3�l.�>��Q|�F|�:;���pD2���/=�瀽ɰli�[��m��k���1�������z�%����h��;h�O�m�hBP�6e�aZgQ'aJz�*�D>�B��4Wh�K�@o]����k�P�|�3��2���Ř��+�i����}*��ca���4��5�>� �ao;,f�<�V���$
��0���>�C�8�y��eROƮa<&�,)�y�m�)���:\�8nb9����# �ǡ���^Ϲo�������A0`T)m&���/A�`�8Y�K���&�#*{��o�����˷�L���L�
���趖n>�|iY�L�1��pײ8�rD<�f+d���eT�cpr,=�8��?�<`��6DF���[.�+�:e!���bBJh��qt��8P?k�%ڴZ�he�$ �N����N^�quq�m�!��>̹:m3�^^�BPG��U4U�[�N I�P�ਲ਼��/�x��NR_ڨ[C"�!2DS���u+����5�_@���Dդ���@mTHY�����x̧}^�s4O:\��.џ�?.c�=	�U%9 ��� ��OY-Ԟ}/�G���s�� ϻ1���+��{h���u�hg�V_,G��v��?;XO*Q׸y%�Uo
���8}�\��;��0JKk�Ԋ�z�����\*�V����h�	d�����Y����vc�V����e��`ql�= �O09�T@6~�T��E�!����?��!����8���ߕ���wש�����(lޟtu	��=��ƍ�PȺj9�Қ��Q��D��X:���������ޚ|�2���Ѯ��YR��l�q̍P@We��=i"�oU�X9�܉���D{R�^8�ǡ-���I�S�W%Z!���/Q���;7�]*�Q�囧I�nD#��[�HO�Q7��4��4�.�:��e���|��d4�3��+�a"�>�6^yusI���^��P<�� �	�g]�3y:�R��Wқ�;��Bz/���u��$���T#�(����Ν�q���zȹ�w��E1��uۧX�kw��|�8�Bu��T!��U��4��mF���0"����^�;�����m9�Q�H�'�uny�����������*#$)e��
��C9ܖmL�?��k�.�0�����e������.$?<����jTR�QK��B�(��UFm�v'.Z�DS�K�FB��Y��c���f�2��t>�3�RaP��0�x���5����!9^R!\5��V��@u����Ol�G�SM���Йo��FL�u��<��(Q
.&g� ���-@na4Ix�bhSGTW�ߠ.�&P�B��]rm�^ʤ�;c�s;="�xt2g������ސV=t4�Cn�l�������LIC;X}���ުvRԜ���kI�yd]@���z�C�C�N[��Y;�����)u��m���h��S����I�.r�Z������ʄ��==آ^�'!��n[��,��V*��P��\���O	E�����O�Ժ���A\��.��a�c��1ƚ�nM���f�����k��9+&,���
��Ӻ���{= [.GM����A��}�����]j���0��T�<��H6�TN+%V���гN���Ӗ�eM5�k������
LsRG�49�r��7�:d�JS��"�H5�[}d?���gq\��W9`+I���8��Fl��cq�g�L-���iW�q
,\x�jM�nD���8W��KWzL�:��pHV�yԈ�]z�m?^�9$Y]�~��ų����#��
g<��Ʃ�M
8��F6�^�k?���/�՞|�N��Ar�����5U"lt�����$#:߸�x����1L���]��t9x��p��	�mB�Ԙ�ibD-_�Q)a��7-xl�L ���A_��6���di�b��l��[Z7��i5a`mĞb 2O�_��"8h{�V�
��
��d���T&���8RaNf��n�V����c�#>��%�q�L6�G�1�R#��o��E��9�o�F��ٳ����.yA��d���,���>����Ġ^fb�(�y�j~+sә��GHl���d�<o��5y�_1W�ja ��F Z��Ζ�8H���`㛖F��E�5~tDcQ���E���Z�X�p麰�����|�V&�f��ƫ�mA|x`��vRL�"�U�=~7=��Fk�Sh{�x�1^�bK`�'o2K���X�4��\��fS'��&�"C�$Xv|҃�O���қ��7B���_m�,�(��q̑/�Y�w��<�����0�����z�W�uB�F ~Q&N� 1h�E�j�������'8�W%>Σ�=��b�d5�1&ӽ���4ȥ򿻘4�Ȟ���(^T�% [�� :\:b�X�/~��"�b�G��;���2l�L*1!��­3j�����#c $yLZ�?E���z+���
�?'cU��ȧ$y���Vl��a���J�c�]�u[g��_E�o�G�"KG�j�!L,�D�W���� �I]�>��Yݬ���|O� ��>%g��?�Z6y�ǙӌS�� <��:�o���kXԲ��a��dz�6/�6�9n^�/W��