XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������LL	��9ѯ�� U"=���w'�5lY�c0���kd\��K��0��> �������[�.љ�rP<'�;=�$?��lQۖ8�RƤt��|�P"��9�EgjV�����"����;UR̸��+����2B(jz��Jr�,UƋeb��DF��gl�>��W��r�O���B8��4�ܢ�&rR\��:-��BQ�wrEg�q���J�� �؋3���-���s��1EWz��p��UF���hX����1I��~�|̲�ܹfo��|H2cm�..ǲm?�t�G�/��.�ߵSfȞ��L�Kc���t�M�ѨՆʘJ���(�Qo��b���{�K4>�i  n��Y�p.D��66��Y���h�q:f'�
�2�n8�(_�����c]ΚV���*�]sD��#OL~�1�����iiĜ����e5�a�R��ON�g�FJ�&��#�K�	"pѦ��6As%%��Í�:�]Pxgx�z�PXGxm(13ߘ�?�Q�}�����u#��u�)~ۙ�����]S80巓�˯Dd&�r6Z�eM�$��׈H��� t�_wED�h՞3���]u���@�dA����!�ӄ4��6��I�2[��9w��s�Z��o6ą�Qf�����ۆ�[�.�?��r��yq��ٮ���9��G��9��N�Y�ǊZ$���?+��Wg�j�ԵOc��>H�Ǘ��j�����=|�ў�!�
�g��l�3T�۶	V��*{�7���<�,B���|�^k$i/XlxVHYEB     e07     680&KX4��}B����S4Ģ�0ՀX�(cm��<���dMI�\k{׮��UI���'��vn���2;Zp��2���t`	�g����va&��(u��C�`e���)��Jo�G�`휹�.�9Go �V��LRo�զ.�E�IF\` ���kwK�S�V�����BВ�2y`Ʋ�_h���u۞*���n�R�j_���:���:�����|��>���&�7#���@�k-�=��$P�j_	���z�6�`��%x�/��X����k
��!�$6o�[V'�lo�o+"��q�gэ��K7�'k����Q��q~2�E�k�P��N����6M/ȟ��c!�f{IMoJ�M��o�H�ЕEd�2�U��E���=q.��J�`�z�ߍ��A�Fi���T��%S���l�U���1���#���S��N��P]%�{�(�����'X[¿e\*�:�\��@̸'o����O���k\�i{D�#x>P�=���~��,⌧B_D<e�R��vW�1>�x�9K] �ꆠJ�PS�~l7��M�����q��ŵ`h!]����~���c�O:SҿX�p���l�m~׊�y�,�A�����W�=*�j�1SZ��]7)��d��+��W���v1�NLmҚ������0"ta�i������@\��l�M�Vd��#�HK���:t�e��"��d�vd���/������!���7��������ʝ���/^��PH�9c�}4����]gL �!��52"Ƶm������#��������Y��2>-,w98&�@��Շ��D3v2m2/�&�F� WR���:�t���xԻa�����h��.ji-���@]՗<D��HD�(�3��*ib���,�kҼ�\�O�b�!Jnz��;�]���[Z��YP��P��MҤ�6����!�~ƻz0�'��B�I5ܗ������}���$��I�{1a�D#�_�m�ۙ�chh�u�Ik[v��E�sɽ�v�y�B���5+kB�G����Vs��;D,w��N2�����R��f�@N� $��G߻�N�D*s\��V. �b�D�xi�&�'��e0�J�탌�����St���R�OY5�ό�ƣE���
9�^]ˢ�q$2>�쑄��.K�$�MfY3���Z�%S�۪���f������#1����?��V+2�h��N��I{$���
~�7�$���X~HP��0M�ϧX����b�P'�l1�����I*�J�_��u��mI����p��r�Z�6����жSL�:��17*݁mw�NS�"��{ї=C5Ń��9(|�]��,3 	���}/S�y���!r����Z|4���A���1LP�_��m>e�i�jbټ%��6+c߀YA���)4X����OO(?K>�nb �;y:�W���5��&C������M�wo�@d�Ư����s`�)c�����2�5����m�q<��|A��D�#�������5zm}O!@jG�.���O:?�h�5L���K6�@N	r�4���PU4EᖛF��ݮCY6��B<vҥP> ;��~U�裡$7���;h� ̾�N��fv�W� �Վ�isq�.�dM��!\����6|E�2�����Q