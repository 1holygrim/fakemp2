XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���G��Z��E�t�X�����?���X���fXnE[�����D�a�����������Ѹ���m�&����C��\O{pVU>��l� ����s��8ܖ��r �܅.����̅��
!wC�$�ѳ|�(����'w�gdc�s��3P�K��S*��*�؂�q��:��؋��G� g����M/W�>{������6��צxx!=�����`�W(ᖦ�%Ӡ���qmz�Ĭ�w������U�	����1�- Wwm��fJ�-&{`G��F��>h���)��#~�U�q	���	6f,F�4E��=>�)$��Bf�]��N6l(83����~����Tŏ==�J#�����(�	��P�s(b��n7	��!�������WW�*P��&��,�R���BC&��gɽA�z)U:�e<��F�#7��XvZ��w\�&XT�&n f	�3�k�f�{O4����91����/�wHp�j����!'B��R�T�7���z���(E�_d�V��-�������ץc�Z�:�ӏ����$�^w%�)TC���@}&�n�Ѝ��	�zó��ߨ@�ۉ0���_|�4@�S�W�X-�-{��0�_X]>J��a��"�1а��\��@lTO�� �ؔݳ��h	e0i�P|l���o�a�0A��ak�2��@@��c�G|��a��܉�@>i�^�.��^��/��,$,�V�P�2��d�>���h��b#����t�� �V�H=س�XlxVHYEB    39de    1170T(veyd.��B��f8�J/G\�n��$���k�\3���.�t�nm���-��k4J����;ż4P:���䬱��^~�|]�:�����h������?�����C�Q#�(���"t���2J�F��d�+��f[�3�����a�c�/b n�x�害BhY3�K������1Ъ���d����}���)Q���S�cv��&��ٶFb [a5R�]�#^�SU@��
�n��)�p)���^��p[`]�[�ǂδ���d���\�9��(��I��},ub����>��|`I��	Ĳ�ޛ�<�[��<�-����-֗Ą�}u;*�CS)V-Ԕ��B��Fy��sZ��$wV8��0%���X�'�;'Px];w&#T>�d��hn��q��}���qʗ��3Z,��.x"�W�k���\",�rG���!u���37]Us)�WH�&%�}@�L��[˷S��&�gޙ�=(����櫫�7{_�P�ff�,�����a�ׄ�!��(��])7���w�H�b?t�@��Ek~+�41�v���F�8sH�RY�5����b�G�vh�)]�=����{&T�]��l���i1,2��Kk���@jcBv����9d%�A����jK����֭�3�>>,�wO� Q���':w��/w��y8��K�؋(��/{���yClˌ�Q��VN!W){�Rz��{���$^�G�3��Ҁ�f�&>��)��=�cG�+e��L���&�e-wr5������i�&�.��^� �odA!�G�<&ݾ���	�~��Q��!HW9{Z��,3%�8��;e��{��Y!uR��z���[^G��M��p�Ȇ�N��C�'�7�[T���^J��e'/uK7�o��" ��{�lP���
*zW0�> e�/�dɿ+�=�8�`$#t9j�����N�~�\Jq�٥T����w8F�>�a\kK�ʯ6������!��,{?mc�@,+Û�U�n4�lIܦ�R#�D�8$1A��.x�C�5}�4���Y�}���Ʉ���B,���%��`��Sݹ]�P��a��������d9���o�/��AJЈ����l��?=j���9�z<���Dц۵<Bf���/K��A�����V��D#���4���m���g���LxÅ�F�}�(�"�x�C�l�������!�9B}MJ-b�zX<|7���.���0�����T};�Vm"�q�c��������?��ٔ�r��2�F����D3� �`;ܰ�`����� \TV�9y ��0�i���C�V̀�s��$��'q�/�������Ĺ~�v��(R����=w{L�t�l���t�x@gq_E����{z�z[�~Dd�L*�x��$�~��c���"�8��%i�MJ�Ϻ��>>"�����L �O5����t(����&+\�ؿ�m�ͪ��xC�����ru�5��f���3@��0�nl r@��2UW��T�r�&o��2S������K�oR�:�r8}�r^�}{���ސ/3�Bh�Ƕ;�:�3��_}%���߅Z�(�����UY����W(�ˡ�`%J�8n��*r��������P��
�5�7%H���
��c���,5tn��P�-4K��%bx�%c^g�~q�x�ua�1���3�{�Ӿ�՛a�[\�
;�g�	���p~7�k{�܏�;��;!Ij��\ܸ��/�}�2�u	k�}^A���}WX�x?[���t������N6��7u�bI��L�{�l��!��a '
��m�F��=�.O�'��������w�X8�?1��.5۔HF,"�a���?�5�j�ݼ���kyI�fz{����8U�bD�� ���[�:���s��Q��o�I]]v}w��V%�d����F��'��Ҏ�"�d�s�w*����{�m�h��z��U=$�� �tZ`��I�	Ң��4&�劳6&�m�*��3iG��Z�Н͹�W�=P�/��"5=�(M��/Cp����O:�0�	�]��v�eq��i��:� ң���>�k�nij���z�Ѐ�n���GE�a�[n�s�7w���|6j�O4V�_z��s���4�4!��g�IM��W���cw�xÁ_[����UPخ�	�c�����#w�M�b&$.L�4紺��z;�����Rҭ"y4"h�E��EnQ⸻�D'g�p)Iк�ߠ`��gd�m@�L�P�+��'��D�rW��Sd倴��Aq�ۄ'~���r����\�R|���-�h�����Z?3���M��!=���J[y�&Q��y5�~Z�)r��#9y�
Wl��b 3*�Qf���7��m��X��*G����'Ó7����Bx����{�/���O�S�Ƥ�~��
��Knr�����_�%��ǈ!^��kĴN���A�IIOR(���"�p%������b�.����A����x9�W��3W�z}�I�3y{�IX�y��wu�4��s��M[�ƌ.�ӗ$"�,��Y�t�taW|i��{�8�TU$ȇ����b@8�S�4S��F�4T�44g�Xev������دΆF��e�z�������S�ԏ �BY������/�b����.��2��>�yLu�ƕ�?1E�~��c�)p+�.vUj?�kl�0�+[]7��O(�ޝmd:����$UBt�y@�Ut"?8��4v���?^���^�\��0.�#;Ҧq���tEK(��i�"�����3�)�l���X��dzU�sTK.�f*��H�:_�'�e`���@��m6c���چ7�Ԝ���<#^*�o]"'DXxO����rB�!e���"�Ya"��Q�b�)5�j�������:���p�(�Θǀ��LX�pj�Oj#���q/_4J �����L�(�۰Ŵ|Ϭ�gK[E�/���l���0��kU�E5�,;Aq�����b!�x�|d�P�.H���4���M��#��4�>,aZ�y�Ƹ��S_����!��M���p�j�E�d���ݻs�ZPX�%�݄��f�x<5o��|U;���e���g��PS�0g5d9�T��xX��Х�7�����A~��"�&��=+Qme$^�Z,�P�U
�P�n�V�)(�M;��'\�T'�m�xF���8@�5�y�gW� �&�,��Oa�`_t',(���Ga�7��Uŉ�s�|�;|�,O�2�ٲ� ����i�^�9�S��$֊�/u�T@�/״��=߁��l�Be3  �G� r�bs����@���JwkE������Y'�T5w��e�x���:����ʻJZ7[4�� X�Ē�;賈��5�2l@w�����1ʫ��I�*��L\Jk}{Ɠ��JbO�Kq@EvX�Z2���ĽVmd��H�0�c�t玽�,Lp0��#9x1�w�;:2B�=ڱ�7#RI�=�,gO���YA�R[��h����Ǜ�N� 2Pl|,����� :���c
��AïJ�o7lp��!���|��^~?�ٶ�	���Q�W9� 	M�赔���MA\���X졎�\���{ �/CJ�H��AK)��bhy hf�h�A�ܞ3���KqC��Yo����nD�����5OY4>��#T�~���7a��Zj��_4�D�������(y�P<k��l�f5���ҧ�ҁ_�&���,�;f��Yȟh�[noWLFi��1��<%��>�\���{j'��z�����"����Z�F{"%�Y��.���(�s�,X�s��������-
�h�*��ޥ��=�NO�`	���y���[�B*�x��w4�Z��'=�Ӕ*�L�aKKZ��ԣ	F��2�3վ��#���m3<����vU�N�s��Zn^_ۊ��ԗY/�0�ī����E���nۊ*���/[��:�&Kw��rؗqy���u��G�I�2ŕ���P`ݟ��_��и'�x!�`��[jP��#O�pCfu�wZ��F���g3O�"+Y�w�8��s�����G���[�T�����}�Wj�6�s�;�U��Q�*3G�v3��g��K�T�k�Ԋ0�� ��Ͱh�}K"y�BN�.E��'��b�u(�(߱��Ï���NOI=��C�fy�1h�iS�-a�.d��8�A�S8ԇ&Ĕ������0 �U�|܋0�����>�z��4�hE�a�4�@��C}�6(ʼ�!��z��K�&��n� ^y=d9	����_K�nDz��<>��R��U��Hra-�aR��Y����a)�尰�}�}Wf�{S�o����$�iW��z}����07rg�!�J�A��^�WLg�^�k�P>�I'��#hԺ�Nvd�U�p����!�B��"(�Z9��h zg�9MNk'�B������+������