XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���X��P���8꙯�����L��j}eӚ2˓:&eM�[w���`����#�C���xM\�._�@��$f�0(z%���\���B�P��XL��\SKR?,m�����B�w����EՃ�����2Ze?[��Ѯ�&�	��F	+��I���l��ʤa���~�ѐ�}.�EYjo��E2N��&EZ��+-���[t��O�2f�����^#^gFub���K�G�l.�l��Vp�j|����q�O�ZV=/���b7�N>5O��&\��#�ֻF'p�d���H�g�о����Bncx��es��]<���i;F��*����#gv�Q��S֝��#����Y�˴'U�y)9̩;(6)N�*V;\��������*��V�4�*~<D���4�&!(��7�t�]�j
���
KL�oR2�pϲY"ٯBc R�'7T�S��h>k�v=9��fO�be��䲨C�Cł1_�e�[0e��To���˱��q����֡�*������B��mT{�GWJ�(:��C�l�R��:g�<���Q�ם�^ �q�������^z m��R�<���y7�6����Y��\	-?��9���7���Ѩ�r}��)��@��K�Ի~sl�C�Zuw%�X�x�#\w��>!��I=�.wZ�{b&t��������j-*�~^���}��$V6w�RK�Ѿ�����[��2����st��F~�lϷ�_P�Ye^�z�����֪L;$~�f
�(���=�YXqXlxVHYEB    1853     810,Z�⠙�Cw/ʻ�� .��hj�{vI�!(ba����)�� ��p�N���jV��2{�%����c;ڄv���O7��.6�a�e �{���O���E�eR�MG��&�s,ñ "9.o歱��6S;5GB�h����J�F����A�����R�@Ȩ�����ڥ����#*y�A.n�LG�oE>i��c|u�[N�rvXw�!��F �es	�#�O�������Bx2�?�d��w[���F%��b������cC>U �u-K��H۠7�������&��:GI�.,t2�m�̼��l�e��͡�>A�A.���-��$u��j��=+���-(��j������n�}A���T�*B������֨������Kv���t� \��f��u�}�z��-}sk�؆�Ą����S<k��
�����v�;(Ge1��N8��������cm@h�����1o���/Ⱥ��/n����h)��:o[/U�c�N�ߡ�/'(�6g�A�9� aU�!�����>|�4�j��>=�Z���mS%6�׹�SQ�����g��R�A8FO����1�Q����Ө!�l�������x�Ȥ�sBw ����M{��MYeU�,�v?�G8�=���E�r1 ��9�`��z��\�2:�r|?��m=Ơȹp�� }��z[(�T6�4gF;IV�Y���$�� ��W�,�� �yh:��)V����)ZeX�L�`�2��-W�x�s�
�Ŀd�Q�f�[�h�D}bJw�*�Op`)�H����6�䎦��ʗz�Z�K��������t�"�z�����0g"Y쳤&H{W�J����KQ'�;�Tt���ʕ�Kr�3�8�sa3g���L`���`#!g0�*o�+N�`�r���NKU��î�M�*�K�M:�V�X�ڀ>Ģ��|a��{�&�̘s�fm�d̡��O7��y���y��)�k���DxL_�b/S�Vr���OD_��>0�	�HB�����+%��?I�
�r�6����y�����*��
!��l�)��<���8�5Q�mtz���=�S��f4>���D$�#��AC߱�A�q�Q��=��,�X3 ��6�Z{�g%��}�$���  񰓪c VF�Wd�&?�WN0)я�-w��Z�>�?=m
-��I��b��֜p����R;
F���'s>F:>n����b]�/͘�����ާUx�M�qw�+��z�r��u�S6Gn�+V�vU���G��]�(���*B|�:�2�s~AJLC�n��Si��k��*ZywVm�p#=�(� �eĘc����Z�+ V4�Yn��=��sc�7) O��Es��7׬@A}�r��|3���_`v��uѬ����-��a��Q��tu�G0u���\n��M��狴�'�毤^~��rp��c�H�\�����M�F��������C��=�[���{�;�	0?a�x�粤Q���9�s����`��W+$�j�tƴ�nc�?��������୞�3��v�J%*%�(9�s�O����bd-2���g�q��X��]�GւyE[k�r���l����ѢO 
qV�nR���`��2P�IG�I=�V�m�w4���ν9����mc�Ryv��}	��t_y����{|��ժ�� ӳ4o��d�����o�V��D"0���o�%���"�$1<�v�d\i���ƺ���!͚@I~s|wL���Ε>�4: �[K{�g��*����mu&]����N/���9�9�q.���?�=�&d�X:���x�&VX�B�ف��;���9�Ė>$ ��v'�L��D��8�o�� z���l���߿\U���yW,�{r�']<����C˳�!(�muچb߂D��ڗ�H-���>���|2�����	>Tb�_~��ȟ���ѝ�U�G�pS�Ӌ��CպKk�����c�"�j4F"a/xvh���8{E�րM���&���a��m���K|ヷx{#��Ѣ��w�8x/��g��i�S��5�$�Q�J-C�>-g��n�{�?W͉>���n[Qu5(�