XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����̄��Ep�S3�3�t���x�%A%�0�#zQf
��x_��Wз��}Q;9ܚ�n�C\��W:�K�V�P�vNH-8��2�^I��i��k�9ϳ���>�c��_Vw�l3�cn�C���U�����q��O��8e�>�K���V܄w��|��@D<$\1�/=(��/��W9V���,�[�)�L*6�Y�9��)oQ�	1[5�\W�qS�6[?8^i��9��Y���j�����)���_W���I������c�տ/H�Hn�T)QvxQ+�I���I:��Tu+���(<� ���2���ˋh�3��Y��W��g2�����K����(F�v��-���� ��Q��!~\Y�)[���5#��Jի��T�o&�����#��C���w��w��3�]�2ͮ2�^C-�Z���KN-��&���Ձ�O��=�����]�+�p�दq�^�F�r���d'����b����+7���@���_��Z��f �XA�����"���f�
֥s�l�1��Cf������+
5��v)5ґ�D���j�8�����T���K����je%��33Og���$#X;�����dqyH#�aU�6LI���L��e���`�oJ����-)��rZg���̬^Nn�i}�������zM��X�!�K�h�Uݖ�Mx�N�k�N4v�md8cenK�F9K���QS�k>x��y9�� u�fْ����wH@-ǍxL���5լ�ť*XlxVHYEB    fa00    2a40o_���0��2�H���Ѳ�[nh�C<{)�w�	��p(�J(T1=�m+�,����[����ʽ�ޫ���(�[�h���}ϼ:GZjלb͖mĀv=��ˈuk�g��3PQ��nT�0�-���&|�_lzT8��J�n���p����W�yt<Ym�z]��%�/No��\���YOE'��B�K#��K@)S�Еr�s���-HҚ���v�" ��;D��xk�/DM'hˌQ��O�j��Ix�
tȁ�c�
�\���nd��Р1�?�}#�䍦�?��2Ɠ�_���(uJ� s��I��ZJ����f4��_G�8 -r���yT��X#��旍�`fzr�q�9''u��������(c���Λ�n��P�f��ې���&�����_��1��}�ycXxvW���S�3���rq2�����DC����>��M&�ZT�G�x&R1[�篓����7u(s� ��^n��g#+�aOfS�K�)��`%"�(g=
p�{���Ǽ"��k7ܣ�A�ʀB4�Hh�yB���EѮ�2��˲���ö6���t���A�P��]���)���z_�4�a�C/y8=Z0��NNn���:����:���ְd`,���`� �e_��_l�?�A��mq��Ņ`T.�q���"��U�D$�oթ�O�!��¶��K6��&�x�LB��LB��)i�]G�$^
�+�'p�X^&>�!�Ðz;�ꞇ*04ɾ�m�)'{��Hߔ�ג�?��͘P$��{�Y3�B�����!���7m���мw'��+aD�F����ZZ3/� 7�e���ܵH�s��8Ф:e��-����c��ȪZ�N�*�Iej��C:���N�H�^z��w�y�ݲ5Q�Ev��93�<X�t�D�NG��CZ��$K%<�h�#�=x,^��fhp����[�����V��ݦQ��l�ŀ��Ū������[c��i���x� 9�$I���3�.۫?�Y����h#�tyM���'�b��cBvl�vb��?����W
|Ɨ:D�ʎ��p����4-���\����ٺ�
YT_Ǳy�y��ӱ���G�gr
b���ή�p	��:�����u�����VfXhԡ�2�܊6b�8�3L������W���0v.w�S:�=��/��g�MQ��4�6�N� &%���(3e��R(`;xq��gD�mW���C��yc��g�	�v�	;o,�O�,�u���ʑ픦	�c;�hi\Yg��g���pE���&�
�B��J�{�l�%�:�g�]ฟ�P��`��P��
0u]��w�u	퉂w�I$���V�,�`�cSUs�ݔՓ�����I~y�r�ƶS�?��z_A�z�׼R���h�Ѩ%�^�"���`NR��\;{0X}��hj\�Ό���Mqm�]�IҀrV��ކ��2�FL��u=уR<�O'��:�".�w��ݮazi��lr��iv�-��5?�ǨYq�0�w�LB�z�Q9��B�c$�O	��ky�p�a;n���0�m����@�V�pMq��Ũ&�F=y���R��VDćJ�k�Q���Q�o�,v�xkC���eGx̆��c��6
S��Cw����\]��X'([�6�*���""����`$M���vb��	�;��� }Òr&��d+��k�����^�����b׮�q�i����ʴ*#�|���ְb^G�)�����f~�� �1hZ�0�_�LH�_Ĥj�&�*���o�,bm��neI�9L�p�uZ?	rQ6��탭�my���AX�n�KE�e"�И����6t\��e�_�C��k�s��:�%l�W��ju��fN
Ɵ�aL���^^���n�D
�7�~��O�ܖ��w���BXI�@���Ӱ߱�.g.C(&�蘍�q�y!��Tek+��Z2���\'�M�F����r�~_�ì��iB{��VOq޴7�ڡ��+I�iLZ#(9_�q��d|
������K��)�����Q��� wP�n~E�@�Lg'�?rE�����:�;�*Dd���e��P;�}R�*��31�S�B����i&X�/�Ofk�h�d��G؆�F*]V���O嬣����Q� L�J�K/�7��!Yb��|��W��1��d�&t�tT|���J�A��u�S@�mx����{&�l4�]���F��R�τ���v㟑���Ҹ(��y`_�N�F�,SR�z<��,d�Df��lz� �W�CR��m<�QS�����4[Q���j���KO#�qWFJ��n@�v٦]s�f~�}f<՞�*3�?���`	zy*7�3>c,̩���v=�"��j	|��g��*�QQS�;�)w�9@��?^^SX�-׿0���19F��9�,g�3�SFx�Z��4y$��+M��7�Jð@�}!��"ہ���}�\ ) y}��)�x.60!�w���H�@?wLT�X�twYǗ��NՓ��{�1�"G��(.�a;p��Sw�?�A$�XC�w� 1 ��f����?�Mn�D�_2$�z�u����g��2�B7rD�z�%�Wz��ѭ���>��hҤ��I��@��;�������0���ut����Մs5!�}��&�(ɮn� uĻM��.N�c����}L_> �4�6�C��Z)b�o�)��L�X{�(�DK��@%͟#��2�\��
��P�ͅ�̰�0 �#�|9e]b<�G��N'�Z��z���5Ѝ.r.펾�҂��Š�Gs�?�vV��T�֪��*b�&�0�!�{� �^<rIC��8> �q�e���)��pOMS5p���~�^����s��>���I�i.>pƲ`=�lB�'���_%��Ve~p�^C�  �A���g�m�d��5/��L0=o�K���{n�n?4�Ǹ�[�d�-n弪�< o���!��ӵf���4G�B�$�y�g��;l'�,}y u����Z�)2R]PĔWԵڍ�W�����������Ȭk�e)Q��X���E~/�<ُ��e>Iq% �$-~��ߖ�)��/|��>����l���X���
����2O�;;N��?��g�>��X��aH��# ��ƀ}>Œ����E�"��^�s������hd:;�]���3,�%3*E[�N>W0����O6�ҷNC��B��Y�F�0]y#P^3yD����|\-�s�bv���,Xˏ!qU񸲬��}����5�{�����ץ'���k8je�*��.6�"̢({�F��m<���~�3�f��؜�1�����]�&}^گ���g��y����>Fp�_g�SzS��ה ԗG~$�Fs!����j)�L '������L'�צ��K|ߨ���4�9+�}ӹ�,�=�Rˤ�<�;rD}ar��"�C|�s�>��o[6T!�����*��;˯��J8@j{�J��c����9�沞 Y�_��ix�~�k�Z�'�Eb��NrD�Ֆ��4�H�/�dZ^�N���N�W�`Թy���9)���u��Rrv�9dR��78���g�0I���г0yu����A�_q��yߝ��}�<����*z>�o���W��g���ڥ(��BF�Y�/D��'\n|�Mt1��Ų
�u��&AC LSc�W�>l�o�l͂f�ݳ����>���B����~8 /�	�)����ϸ�ŇFo��/L��'�����hK�yߩ]8��0��^֛ �v�i�t�"b��}�����z1���{��h�r\��`q7N'��u�N����\}4�|`&`���HN��(ޕ�T�;f�b��5���<����>�k�!Q�uT\��"���h�Г� ��؏`�5E2����}�_ܚ���y�s���zХ����[�����ӾO����Q�H
KSm\)��9d^9|.u�h���S��(��!���P�lu��c�:ZU�}g7nbEɜv��/a��&�����Ga��'7g�¯"�C�=K#�*�h7�Ш�)'6O*��ۚQq}��2\("{��'��j扢	$���g��r��*�ƞw�ٻB��:.R>�<���L�vum�<�i�v�{� ט������me)\?D/56�Ϗw��Y�>B���b��t��.x��c��>eT� c�F�,�Q+ݬ�ѿ��^����]C��+�����~�����*o%��x�h9R^O�DZ~�[���1�o}#]ikɃ\%*�h�!��9ZAѷ��U׎��&�O�x�D8�V������Xr�%\��M��ҝ/<1��N��xT_��f_�qǊ���Y�ë_�ڳ�	��=`r�r�J������ i�r	1�-�Z��ѭ���w�խ��x*Q=�a9�i�R�̫��8_!���.x���|̝r�~�mI^������[��[pcqP*�h@5��r',6^3>�ML�qClK��3\�� 0��i@!8��r ��PՑv�q9��(D�I���ծE}��u�$ssa���>f�3�jJ��0�b��y�pp In�hh59oGA��c\:�R�Y����E��_� S�e������~��9,�`1�C�������t�Tm��Z1l�o8���Yj1"��4A��b��G���љۚQ�k׏��X1�V�cD��G�����D�5M:�F��н6��+�xP@ˑr�~yѵ�pW_��1c��#�@s$8t�7[P�'�ul�R`UJ��4O�V�2!�S�5=ܯ�\2���Ɋ� k��0��k��s��
6͒�FfZe�1���ʍZE�ؓ��Wt?7�H��l���'��vr������u]�e���[�S�r���LǱ������H���EЂ��xz�C_���/1$����B�3lJ�k�����6%t���Ni��D����v���Y��Rh�UF��j��.}�I>��X!��~��]�~��^y�ld��&�?y!/~� @�˸m@:!H0�����g)�X�g�j[n0��V���-hiؓ$��L�.�tm�Շ3�G9��`0K���j���A,�}zΓ,pAB(rd���X�a5��r��y��[2�h<^dV5e"�[@���p�V^Ef��
�
��L�?�g/^�]|묹u9(I3m�s��̨�� $b�n@p����2B/�^��+������# � �g{��k*�;Tݢ�8�I�Ps�!�ϔ.BlC�ψ����v0�����:]#�b�c~�7����x0w�c��V�VB1�Jt�\zEu*�ih� ����N���HM/���1�`����ǓW䬎��r��@�R��Dz\�YՊ4��D���X�a��KC��O���Xa5$f�`|�zfG>��H��~�MF�|�dK��L-��Jf�������rhn^�$tKі@�*�������f	q�x�aߏ��G��OTI�Xw5��]tX�m�sK�;i�N�i�k1�K�d��*A0<��c���5�I`+����j(|���b,�D�5����BZ!��Ւ��Jn�_�GN^�6���{�6c���D:],dɼ�k<`��35bO��^C��Q�g��w��ɧ�Us[�F���R*E�@C�n��S�ϻk�X��mS�0z��8�rjx_�_GO��"����L��4I�SkC�*A(g�Qn@p��i�'L |巘�En,��x��A
����zd���2��G��t�k�'?6N�5&F�▍+#k�:(|=�T�(�i��S������;m���c��S�����7Y�����ˠJ�-U�Y�%���W����3�A_� �9��"��T��`|<�a�毒�����E?H� �f� ���䜒�_���.y3��N[�o¼�]�vu�H���e�s؆�й�ڥ���m=����E������1i���)�p-t�+����&���(��ǌ��G�ZN�B���_':gR�a�ⱛ��d�3h��PwXq�v�*;l+)�� ��c��*�mf'W��A�@�.���?����[������|j�������hB<�IВA����ℕ�S�������%��w!\;�l�	�^�w�~���se�P�D0}�Qs5�U��Cx��a&'��9�ɦ$͹_(��,�s�*毾�ը��*�*�ld65ZNK��b)��2�}�(Q˼��Mi~_K�B���N>�|t�3��F�1c�� F5겻��z]nf���B!�ͳy��K�-�����-�hÒ#$���]}�E�͂{�b[���H�&>�štr&vY�XQ�0!�0w��g>��bذa$dvoBĕ�}J��Қ�I��uYd���+\���"w���GĜ���O�|�p�P��=�]U*�t�h�k��-R����Z��)��%���߼���=���s�겴�Pey�^+�10�+��,+�ڳ혻!�=C�d�s�Nr��x�vC�O#�3�0����o�f��INk��Ѹ�oE��HL��0伥X͌8����7>l�������W�~�K'��)2�O�1�1?����pֽ+�@�8���e%=��r����ލ����+7���=���M����DW.���q��85��y��1$<YR��l����i}�w�ڜS���D����U%����Z�Y��Mk���B[eGX��;�M�F@������G�y�䒋uZ��t�lz��a0����F;�8/꽹�}������K�3�ؘ�%�6��}�`˳P&3k����&�V�1*�x��?e�$v��v�1��cHK��m�R�l �k��Z�?���7�V�6@8���Dt��נ�{%�Ҟ��f6��a�Y�O�|	w �,�=4�n;�m�L��<�e�e�ƋG��wX6�O`�4E��)��� �i/ c�^P���l������z�-D��楞w|���A��u���w�����-�20��Լ���!���lc��V�Y�-격$ �m\�>Y<����Vk���5�	�������c�x��X��ٚ׷�3��H��>U�k�M	��-y�-�{�a
lF��[i�}��O��_ EU�#�ؼǐ(���?帲�C��Q$���l D3d���N}�-�i��h�1N&��� ���4V��0f$��P�o��+�!�qS����Y�7mr�3w�l�yojT�V�5lc>gGK�䷳��́�9�*�A�k@��J�N��9	�8�|Ƽ%)���*ȧ��s5>�QI�NoED1wl���A�t�l�.���T�-F��2�4���5=����: Q4��s|��/�-
��@��2:�������R������{�L�ЕKt|��R�8��Z���A�4�Q���M��M"mn��¨X;�
e��8��1M�S\G�T�Y$Ii�8�n��s��
��~������ʯ����P�e.�!�q�q����y.���=7+�:�\��k�b�{��
���y�c/h{� B����h&\�/���Frޏ��j�n���u��nVK���/i��3�0Ԡ$�3�M�Wf���u�$π�E�����ф���C��jgGc%�F�Uʍ^cZ�mqYA� "��S����P+��U���#��8��;�������+�)�D`�ܛ���[V&$4��`Y��
�Y������*�wi��=g:/
����d3"�+{?�����V����_`��9U:_*��X%'؉%5af�Y�w�;S<��*�4���*���������$U�1)�'vJ�f�z*8� �7���A3R� @��=S75�.|�F�P�U�ڳ`�`a:���9��{b쿼̻%4���;I�e3����9'�Rn>������뿚9�"��y��WA�I;��&�O����M> \p)����-��TB���h�]����{eh��L�^4��wf���u��mi���3�Fj��E�nX5�x��[��_dq��+���8W����U��p7�9�
�	b�)ҭ5տ�6pA:����peHK{�ыe'J��k�K�!�0M�m`v�iW�q��!G|�!O�U�Du�f��L�>^J7�Y�(��9��>��b�� �-�����@���1ezȲ
���L���Y��	�<�Ϡ��������#F-�/H�.>�����͓�;�\��ǵu��>(Q�ԋ��(��5R�]K@�2�1�@��<:v�V�f�z�G;���eW�D�=nB�kOE�1��"t��L�?�H��SAGV*��\H���X�'�
�*CÈ�����4B����!}h\�/��ł��!|��f�Oޅڧ�3�pl����!M������T��-{��s�\�C��F�&[/"W�z�=���փw��l�V�y�1��%�y�N!�a����_e�|�9v�9EBЍX���	e;0Bj*�LcA��m���S��p��UY:��Z��.�S%��(��[�"� #ޱ��J��<d�d������{��7�}�K|���\�)�VJv�]�G�x4N�ҴW�V�9x[0A��`T������W����D8m�ƂY}з�/S,ߴt)�V����ʶ)�=E�{N��H������
ʫ���vF��C�e�n8�w-���旑f�>+19AD�R�^$"�[c�K��e�&湚��������dN�?� ���/�}��Ě|2+J<�4�"��!֊Ŀ��:��6H��{w�'�����t�T
���+�A����Q�����gʏ����>�x�I�-�I����π�QG~p)�"3�`p��!O� ����o��,�*���no�o��>0���2�}G�y7�z�;�6>�x&�
��I:�Le��V��4�GF�Hi�*ȁCc�|3�����p�B̓6l��҃�1�a�D����wgX����'���T���L'\��l�CL�7аʯ�&�i����8��LJm��8��ߡw����*U£@�Ewl�H���Z��	�paF@y�T>�Y:�5!dYX���G�͜3�;�0>��J��Aj�]%VJ�̮�^	0�X!Ex��w��u_:�@�mF��xm��}
Р@�$*Q�r�F��@�C퍟I<L��W	m��*��: ����h���k�l��.FE�&�L��fםG�; S�]�p�� I�lػ�o�(�%M��. �3=���p"���ٻ�b�ʌL�D��%�o���Ki
�1wm���(�]"s:Q'�)��K�<r���{m�W���+��=ݹS���%�m�M��+������g��驘}V[������]�Q>L����ܖs���"���ĆĒ�Y�̣�=��2<�/�kd���"JAZ~#����d=e�e�ʌ������:���ҡ*pʟ�� ;��rU�bd���SV�/U-:��;�ڈ�S;�*�2!��p�Z(���H#�i�n�%��^ԫ�]۫k|��ό���~�����;���|Ѭ�iq=2�Z��������� 8W%Ȋxo.�?!�͐+Ԫ�߷�i�� 
?�R]z��I�x�P��,��+�P�9D���$`^�����h�焾�s7 4η�Ǡ�G����r^3�P������o��-+�\�����w���Bu��`A8��Q��})Ab㈍�,@O��O�Gul��V-����O��;�~��Z��t2~�^�1c�������e$5O*H>���סk�8�%��A�sY�x�~Q��h�o&б{x���yЃ�� ��U4��W�&��@z>�("xe���0�j뵏�_u0��DX�� ��֠;��)Wh=��������A\��a�$jc)��/,����g0��2%�M�=k}f��`|� *5kl$�ԤiYѡ������}�	+�Z����(��k�����F2��B?Ӽ�C�$�{-5?-��ϡ�Y�e�Y
��\�D�g�!��q|�Afbw'=%1�ٕI�	Y�*�f���_��C\�����fgq��!]M�̰0���T� �-)�,'�1I�����%2�l �<�B9���4n��?�|����j����"F$�C̎.괴*r����^i�7�,O'�U\��Hǒ��4$�y,lݝ9A=�(
���T	m���ӌ3w��r�@��&� ��GW���0�a
h4#Q�����偠
bJ�<�T�窼��Ԃ�8��������E���^�e��6)�kt5�~��0g��I�hs �MqޅdA!��tT"Jm�5��Y��m�D�5����I&��Ĝ��F������ xN.jX��{J?�?�Q��{ګ[*=G�a��M��A�;�9Qlf����D���=�z���}�&{6dϘ���?�Q*��s��d�Rl�EiT|>�ZPbO_ȫHf	*ަ����!�hM��X��y��ԟb�� n~�����m�����f����yZ�y�B�l<&(�Sե �U  [��eʱX���l��S��Tl�r�(8�7�B���y7B��#���%x�\�F�f�*rB.�Tr�5@û�C��ez�m6y�	�+��%*�+����)�ƍ�H�Z��=ZT�����f�jv�qL`"C��AB��$SԒ^f!���Ov��g�m�W$��؍��*ʻ�zKU-��F�M�ց�}�
���.V�͸��Sh+�Ǌ}-TBc���o#��Ҭ�o��A$�v-0�e�3�� �z���k���5|
�R=���$-��Q�ɀ�������n=.�/ T�U��P�,��4oIs͐�]n�Sv`i@�Qs/S�'��S�O�ىE�
|φK�mYPkh5Z5XlxVHYEB    fa00     8e0 w���[N�X�t�u��j2��~�`�����8���i�z���p<}t��},lۛF�����RW�ώ\9Z�l¾;��w�;��8���$UX��L!��P��|҃�.ļN*Jg�$�Ns�F�/��¶,���l?��CU��7�W��^x�D]
����	?ɤa�yY�$^^�x�с�כ�Ϸ!œ^��,���r	��)�GD�T�
��j�����o|@��\�:�����8��/>Oq#��T'4��X�r����G!~;�h�3����<ְц����bB����v-�eN�����c���Q�}�䰋�n�1�z���l���Nx�B6��χ����E�C
�V���4N���sHN�ڣ	6h{m*�rFh��>��hgV�-�Ԙ]z���e��N����DkTe�ka�����)RvC�w�m �ޝ,��B �@��dX\q��8+����`�-�<�)�Qh@����:X�,4�ぢ�!�͔��/m� �������j,�gk��Ǯ
����2c�+��Y�#��I�Q6e��6r��HA��Q@QN�՛ZC�bhю�z"�|������.�8 ӀB�u��X�c���"d��Y�B,'>��G�b����!o
[m���)����Vxt�"���$զb �OH�P}
{*.~8շ0�o�hT*r;0O�*��O4Q6``�~�J�o�թqo
���*���!�i>�Yyz� �ީ~؄��;�y��XC?h�mA&E��6(%Dl>��S���m�\�4�&�)��Q�ㆣ��A������S��3.[�*���5c�ŋ���:L��9AjC'?�T�>�SO������3������}�O]��K���T�r�����<������k��Z���2@��n�"�������j�j�!о�F��w	�m��R��$�����O�5_��&�tg��	��#r#�t�?�5.'g���v��k�O8�Ӡ�Ӷt4����_��Z����� j����3ib~��Z�{���[C��d��
��l
5@=W��b���m?������2Cgd��cx]�H�o�M�Ј��%1���C(��۹��|R1���z˦�ܥ���Rž5��*:�q�N�sxv���7��~���Yo�%h������ʠ�t�3hD:?��.m�Ѷ�E���r�T����������� t����L�����
{9%�?i�@T���6�s yJL��TO����s����	��x��$OW�����S�k�}͍�|�ŭ��1<��E�I�ٿ�J�l�< ��ƍ4��������$�����|��;��^ @�Ur��-�F��d��=�dM���
�G(��P��'��Q�U�[��7��Yɭ��Yo��I]_#�t�N{�z:��}D:�0Y�sz�k�-��HЪ̍in��r�u\��nV.�Dlh�L��?@����_��y���Ćg�zbM^��i��w�Ӱ�q�X��dk�[3>��׌p"��͎�ȋ����I�}�Q�[ؕym8���`�"9�o�� ��c��X�,�Z.*��٤S�݅
_ ;	� ;s2��M�i�0��?|��%�>��H#��t��8��n��p^0x:��&�FZ��[����͖�[��]���.���|��α7m �'P���X�c*��[�1��;��!�0ʷ�����e�]7z�J�#��:��lb�f�\ֽV�(?�޲t
��MF���D��ҐU�ˮ`	�)G)ո���x�#r��+��,ͮo@����@aۃ��C>�b�[�J�<�M)�:��*qǝ��_ $�	-��s�N��x`:�`[O�P �CPl֚~�7���٣IS{ gsL`(�=)+�X����*�>��]�m����0�-��>"(�c�A��d�gaMc0��{�2b	�Jϰ�:;�V�Avux��:3�O͑D����n��f��;����?����[r�3T�B�Z��2e�5���Sj�ɂGAs�Ԑ�#�p��8��l�1g�'@g��Q����U���%u�J+H���l�G�iޠb��i,��n��6���@�ګ���\?��.���$X�»�U�@��U�)��M��\������uN�{|W�x�+�`��� 7���A�R�w��>��`a��Āf�u' D�h��G�.K�j*�{]Ӈ����-����f�]�����Ő���A>��`XlxVHYEB    fa00    1110��٭X��S�_n"�{��xz4��nO�q643o�C�$Uf�w���Jx�9cơ�#yҡN4}���g�e~�dm���P�����줜R/o���O�����Ŝ�_7����7Qw3h�}�?X�q�S�}6q�K^Z��p�;�!���c�!F1�W�Q��i�r�.�8���L���8�[����is|ݿ 8�}�76�	�A1VSؤ&�Ҩ6&D��	�=�P�v�� -T-u�n�4��6�%q>��M!�+�5QK����V^���(�?�R�x���3��e�Z1Ik-�3���/��^%��,�Q(��TwAe����0����2[���s���p*ń0��?#>k�Nt�_h�ız��6�&�]�[��*[)f�慓6~Xy�q�����=I�����5?�e��R33dAƑ^�}c����0)>�q+0r�k�X��^z��J)d������O���ꇧ�ӄ��S�s�? B���l�
���֮��ԩ����N~8���ݻ*��M�\���͓8����׹ǁ*$)�n֚�(.��q%����`^��JK�u���Ϻŷ�[+
:��fʨ��${w�f��Z2����sS
ݮ}"l/�bJ���R_��R��s��(w|J>��-���v6!�Ӧ����>u�|�>��~�e?5�:��5�N�W��f  <*�6�C���E�ǜ������Bs�ڶ�f���O�C������;A�Uњ���M�R�Ђ���⮖ۨ�	�]��*~n�E�m�=�<Gsq+_U*a�`��F� �;>n�ԝu�q,�6_%�DE�1��� '9{�1��t�,��i�i���,��j8~n�[_U����5�������"��g�a��F���G��b�T\'�����a�f���~��$&nȼ�^�<��鰓����pa�d���JI}��.�s�9��蕾��͐��"H�	m����WD΄�б��]\�s��[�I]^�̛��D���%pz}y(���\_���5�j�V� [��96��]Ι:�S9����A���߄m�5�nЎ�=��X��+y�mF�j&j���Ǐ�[��H�7n�h~»��𸑝V��}B�-��R�F?�8�Y@ībC�p@nin�(���b0a�Yh���w�_�.
���tZ9D�t$B)�5a0�J����
������ׄo�b�mUpu�,짉�a��:�˾</ͿHqn����X�O��T�FDU_��8�S!�����DW]���+�76�9޼KC��G=aV�p2}��U$�"�uQOt2��6�'���>Ȼr����Wc�,P�
�������&���O�K��9�.(C�B��'�\	�ɐA��6\��r��?�WS������n���5:u"+|��;�Z���u$t��t߿�"������B<&�C�����3��7 �y�A\|=ɦq:34"@#[|>d�OYk���o����NҀ`��y�f�vo�`���v�֮$�8�1Ux��AK�Ǭg�s_���H��&����P����z@�jfo�����*4��,/�#�&3� �	�C>>6��S������x<�"�nMCh�y"(�,����~��.}�,�؎�)��s	 1�l3rS�6��PQ#�5�(C��$y�(s��Ϡ�5C�-x���Y� Pd�`	[�ݥx��e�%I��҉x�����T�������w��RB�N����qG�#
h�lԕ-�U,��U7�Am|*��!���m��`��`�K|~p�5���V��J���g�?R1;�C/�'v����L:e+������9����4|>/���M@pU����r���d᭜��A�żA�ѥ�r����X*{n!�������Dx%���]��=:�+���h���1b��8��GO�/n��N����8[��L��Z��Ps��8�߮�u���u�M��-K:N[(uʦ�9�}c��L�v\�q>�4R�q�~n^oʇ�u[�]ǊŪ)�\��?��r�"�6��wn�7y*u�a�&��5�� M�Dvxb�� F�f����r6�C�nD������t0~�7�Ț���;�}d��(\N_6�-Ha7���|�<$gB���y�,�A�������X/Ϙ?�R����A������T��
Em%��,B��$4V�0�n���k�p�F����餤x�!#��S*�Û������h
�HJ��XGrc`c3�N��S�bro��FF�sauǅN����p�I{#�tw�]������EŞ�������Rq�C�v
m�5�E}ku��&ǟa=��e|�$��L�j�%D�az$����/��+���H�|+�cV@B��M��� �J����2��2���o�t�7����e� 2�0uj�רY��o�>���l��\��/��p=::�!�����F�����a"���Ӎ�ȓp���[T�ȫ+�?�q������Uzy��~]Q�e���I��^��_��R�����_�$9�}�:�'i�Q�p��o�^���Xb�
�K���[�Uޱ��T���W��R�Z�_�x�_�$� �H�1�8Gư(���%�]:(�0x�)XY��ă�8hv�E3�H)���y��K�SsO��� 72���>}7�`��!ra��Rn�^͖��6�ӣ�<��;}W#��}hlo%�1�

��/��Jhö�$�'yI��~ T����1��oV���,+�Di��:�s���|�����ے�ON?�`���K.�oI��+�(�g&��eX��­���G$�܆�ȂY�e��`��m{}�����s� ky����4�m� ���®�Dv'}h>FK)GFLD1;��QA!`��0r�y`Q0�b�U�MGuq��p�%\�v�,v��a��@yU���L�	�*x�7Υ���`��Y���4޶����ܕ�8�\�d<
��H�3�f='~� �ov��N�|~uJuj{�1]�L��Y�ͽ{4����׼M����'�	:�f���#�R�W�(�"�pI��f@.�����&����3�c�W�|�g=�_�6T�E݃oV���}�[a��Je�S�����z�Md�	�'l���N���x��eg�47����D�s�\������]#zS�i�JE��K��o8ե,��,l29(�-�&���w{���t��6���~:�1����mtSF_��(�J]��F�}��LE|5���ͷz�`I�|ϐ?��<��yv��5���Qt18�� �Lǟ[�2�.�<����1=��kŠ}"ؙu6ġ��c~`�Xk5��/��o��q�I������C�����$�&A���L�~�-���8���CO�?�P	Bz#��6��!>R�1�OT���"��&cE�lCn�c?8ȴC\�O��F��(�ڷjצO�2P���^[f=j�F7��~��u|Pob򓅓4����+�^�F����0�X�Qm�J\�6#b�_�Jp���"��Ũ���ŸnH��,���UY���lexL1��������-�KY���*���:���Й(v��:�s$NS�����q`����Z������ς)�G&/ ��'��ߕ�L��T���!C?���9Y�HYce�����Y��-%�e����O߿�e�3� vρt_9���.z�Z[�1��� qt	|?w:u`'�v��'�5 t��[��n�.�PxЕ��+M���y��@�;!a�~��W��f��T-�ދ�9Wa�roLc�{�{�7�`����?K�u~�EOq'�>��c��-%��Ǹ�ΰ&��v}D�),�ap���Ͼ��)�q�Z	�1��ӣk`��6�UȁL^l_I)�u{,�V�tI����A�T��	(�U��mNqFS�j�0c 3.�?��Ϭ�����gm$)�.���G�x��Ee�k��y�����-��_!X��n��#wj��/�^ ׳ָsao`�I^T��2!W~�0��f`�,
j��vV�!і�����5���	Oܡ������L�;�-wN�`��2�M�1��	��@�p�P�+0�+(�(їr�V���⥰�<=G���'�F�I���2.����3Z�O���f.��Ǔ��am����-�ƆV��A�+K��Fa���slM�^��3>*N><�`��(]IE��G,�b$����\���<�봐j��X�솭���63c����������>W.M܄�/9&A_�&
�l�ӝ_���ޡŲ��l��"�^_>�fc���Ւ��Y�=�/9?�yF5�Y;����+[�=ȳ��Ҍ9J�\RXlxVHYEB    fa00     ca0;��פ�j��W������bY��P*�Q���0������Xc{�Z
���._o�3ֆFB�t�B&��Ab�
�q�p���O�Uu���Se�mL�W��l�7Gt�-��jʰHQ([�{��G2���ɆM ��*Fޏ� ~�j�C�� �d_��-�B�o2Q��0�ը��*��Ϻ!���_���Å?z+��7:��'ž����󺮒����#��Wh��� �'Z/iL�̯�z��2�Z�a1��ݶ��2��2 ۤU��i����k3WQ�8L���=�u�"W���8�Y6��	L�{8H]e ��T�vc����FK�D0�5�-<J�S�X��c��U��X�T����Z�N�T;(����{�I�)��NA�RXkY�����n�:�	ƚ�$��ndх���: ��{�Zs!���i�09x�9�Eǒ��i'��~XU ���E� Z��A�A~���j�E�����g�S�恷t�M��"m�L�����N\m��(λ�42�D�GM&���o���n�}���#���;{�)��CQ�X:�Z�o����L�������OclE��(�h��#��i햛�؉��Yp�=�	 ��2������3�nQ��6 ��:f"n'��F�^W��`PgNPDy��
ցT ����7H����fD�J��yWj@�{�k)0Z'-���:M�MYy���m!��wZ���|Ѓ�J����^e��&H�qr���7;02vZk���y}�g�uL��TSo�p��w��c0�f�E�e5'��p>�������̜:#1�o��.g s?\��=�oj&W3|F ����]��>+��}�<A�su:�k�v�L�`+��Pp��W.��[S�!+�>����N5A�/ab6�x��K<m7d���p�e�x��V�X���U��Q��f,ٗT	;��/��8j������a4*�m�q����nY�J��-����g����'�&����A:Tt|>4�v�*ۢ�&K��qMIT�+O7G�C��^���]�gPq��!�Y�����F�k.C��M���S��w1��7����E;\�IM�ǏE�q
�� ,mc�
sD����Nxt7����Ab�%9 2LA�����fs;$�t�]j�1Ao���o�]@o�}�El�cDθ�(���R
�X23��d3��~�r'C(���J�6��[������d�%7D��-��Q��kT�j�zW�)B��i՜��Nh���d\ѧ��V���+\����o׿i��ʂ��˫F�ݧ�o���}{�;�m�q�;H T&
E΅�� ���F�����4pa}Y�~�#J���\.�-�Sl��P����Z�șv�rѤ-��^��$O�]-y(n)Ə��A�3S4v�ߌ$�~{/������L��h����Q%(�a���9�c����a��|n�A�R�l����bÙNaa�4��+�O���j�h�2�<��ר{��,h���D�
.Hi�Χ��z/�aA�#����ָ��DX��Y.r?����}���2�?����%�]R$6��Xi�5"W�`��#[��W��f�����y����
0��A�d4�2�_�|��Mn
���z��0��b��<ṉN��y��;di�h�Vx*=ұs�.������6�b���S���T��j}W�_\0L�������n��|��cK���yu��Y(Iǆ�Y���d8s�S+򸘬�7����R�h�Q��i�K�K�F�����1���b~��%���F������YF�� �#ػ����Py2�䨏5S�1C5�c�2�Ӳ:bۻu;A&��nA2�J��!t��ir�u���MMƁ$ΥՅH��¼�%�I+��O�l���.��IY���ԣ��Ӆ�rڏw�5^iU����3 ����m��?�)Z���X��'�ppN�-�Q�6��p̈́Դ�� .�jm ���.]�[vNT�3�4ђT��/����� +��p�N3tR����3��{+�)�����᥉��t���Y�h�{����鄳����B�d�a 'ӿ{..����N@gmD|ne���MvK��a�ɾ�_�=|k�,øn�u��U%S��� �?����8�G�����*�7;���/'�;�}�4������WO�F�d֏B��ǘϰ�u��hh��.��>��d�(�emw`1�ECX��~&º� Nl�<J(�F�*�qs߃	��@��%�],Sg���$�^�:��?���q�c�����?�.M�:�����m'�ËZCI*�4~/��� �[�����}YA1xo]Ď#�X��m9�:8�g���uHl�mrZ�09@Y>)5G�zB҆=V,��@Ĩ���c�Kf\���G���S�]�#�c���lmfb����H^6E��n S�qnu�06��O|C�` H�]�b�x���~�v�q�S��x��>#�ȫ#d ���) �b�����}]�nl��ś���l?9��� ���8 Eix�̨� ��ՠa�[�.��oW�����7�{.s�(R�m�G9�٘�`yW��㧁N��=��/�)�$f5�5
^\�����U[r/j�.8�r�䆨f\5�k�C�5�E��z���dG�����E�qWw?=�l"���`c�ɰWZB���/C����J�ݔ���0t$�p�l����
{d�Y���4��w�$"�gU(0`�$��
��s���6���"������~�iWgY-�[�'�
�I�6����'>�]غH^�v����h;^'�I
c��!Y�KY����KkA���H����?ߋ�ħY�*��p�����a��ݶ�jt��J�ҙ�F��|Y�S&����T,1j۽��F�n��d̊`�%��Xx�lx������,��@������67@�P)������k+')тa�"#l�^Gd^b#_����{�A�l�%D�G��e��!��[��c�%��=7��W'n-&����Zq��k�+�;�T�!�=�K�(#�>���?3%�0���� *�9�s�ܴ-N���{����|��LsP ��HX��)~3�BD�
��x'6(��#�,��( +;S�-���i�����&�;� Ê�y����N��s�ێ���{)Ζ��
�c��XlxVHYEB    fa00     3f0c��Ҕ��l!s���c�<�%�Pr��az�"�pb@�Q��s=������/�>[nP�V����`U�:5O�~U�A� ��0��U��P���!O�r濘j�1k�ȸ���S�5��h Ԁ�D���%Ɠ��^��Bv�V��<��B5P	���\�M\�X�0�Ē+O�d<�v�G��/[�(�F=#�QCA<͋ �"Ӈ��W��̋��A�7m��L�ɾ"�Do��ĥ0@�|m�מ*��<ՙ��R�q@�Z	-H��D��B�@߂>�'`���s2�͚�Q"������M_�Q���;�]�d2F0�v�0�b�Mq�1
Ŏ��Ǡ��y���:ƀ �G�eh�
����m���/��g�0B�-+���U��r�~�n��(G�F0�ş�7�ߧ���:����m���,�1n�??����`֨���8�pq7}e�ߧ�듗�<�����%\6���ؘc\���� ���X�p�-D�����ח��V�?L%x=x-���;�>���ȡ�&@��t���q#@�R',�N�C��[,�{����_Ey#H�Tw��Ll�8*E�̴�O���`J�pb(;�Gvˀ4���Z�@im0�T>~S�L���8����gy�:<�XכL��?�щ��.un��h��y�7����w�Ű�B�r�+1�U�z>�f�^֔��IT�n����9�jGߎ,�5�=M�k��[!ه@�s9�Z�t���s�}�s9�-�$�-��d���6�)��0�F�R�ҹ(��h�҇�q��7���A��7wZg�o��]jUH��x�M�>7^�밃8�;Ż��x���I8+c��A4�W�v�7<ں�/ӌ)@��(�Zq@y�I��i)� ���ݣ��:���VU��w�V���C��6u0�j��$�skiا��SM����:��ű#1��?��x�q��<k�ݝ�c�o)n��1_`��)-�вi�����+��j>�5o@�<J��;�6sW��v�,2��>o��c�	��XlxVHYEB    8096     b20�t��vM!bo�Lx�!O��y/��n�񤜽ǲ������o�D�d�wQ͈. LBF�`Aۅ ����]��ѱme��]�&#�VD�@�!�g��^+Z�+�u���s�l�By�,	gna��5X��1T��=
�G�O���P�O�}�6+>
�
`h��E�t@�ΔŁM�7���nC4���[��%���t��,���Bl��(>7 7�/�d�1!<y������;��Y�N2٫�!.�lRik��+�|�%R������K�\������BТp��^3������]���CI��%oj�<B�H�� �
gQs���5��yl���1~wg�כ���3��qe�Ic����q1f"
,@�E�2��:��̙u�
\�nͩ˒��Լ����đ��o�{9�׀7��,?Ύ�����wɞff�����'���u�����Q�U�0�T�ǜ����#D%=NGR��<�K�QO�N_�@^f�������Ov��{x-36�$�����P��N�H�G������b���7E#�*HX#g� � �r����D��|��$�~����t�N���9���L>K9[Κ�.;]Q2�J�����Wm�V��,��-�9�Fޜ�\ZZY�|ׇ^p$�&Kf���n.�V�9�B._%x�?U�j�3�s�t�����ƃ�ޛ��	J��K�oۡX��Z�9���줰cN�t|�uQ���!��hiK�x*eq���h�L�I;f�5K_܈1@O�q�o�
�ZgS3��h�~����;2��FaIQP�f?�,.�O(Oɨ�G��nӇ���6z�Wv�L9�VF����.ҲUt���l�V±��j��7�d�ry3��$U����{m�6³O����3��Ӟk����?<7q�� Z�C�����F��c��4�����I����4�u>|
pH��Ѥ�b�z3s��
�?1��Rʹ�J�4����M�$��y�.L�a�B5�+�q���F#��,��m.���ٓ�,��t	�<��� 7� >�5���#�0(O_]�G�-��Tm��\}:T>��svU�<�$�D�u��[��v����Ly�ڀA?.hP�4�fE�+�X�Č�F+��Z@*ɮ͙`�!��s��_��="m�d>�S��HL�\Դ�A[�jl`��tB�RD!F�87Ps].�G^���<Z��rM*��Xa�I.�: 0�cS��q�"��f_y&�{;�m��p;�����.8LK��$�lߓ���^b�&��U�v=����|�]�>o������d��{)8�"��D-u�z���,�$)��'?���R���\df��RTo #e��uI�5��z���S��3Of J�N;�0.l�k{��87�����F��l0q���pq�����m4i%�;��PQ���{��<IpTV߬$�͕�q���P��p��V�G/���kX���u4l^JM���[:�k�m��©2�V^<�Q��dH\���C�{�0�6ǽ3jP���![\jO��ηs�n�X4bڢ�i!eLG���E;�?��&	BQe�o��$寺f���������
��^fQ
J�S	:�#	5˙�x0�*�Q|dԚ�~V��J��:̦{��f�6�}�:��ә�l�e�7.5|�A�3עm�NT ��p������L]@�pH׮�1|]��nw���P<p���7վ&v 8ja�LK+С��0��q��¸V'(@g/���o�¨�"\䓓�	�M�n�#GC�49�k��`�.��)�8K1iIg�k��������/�LU �W֢�o�!J��x�
e.j�i��C �z��B!�怄��(z��@M�ja���gur���m9���� *�Bƕ�+�h������}dQt@U��B�kn����!5+WͭM�(����(E�p�A�9+�7ła�?�CIH���N��:�V�p��*�r�Q��Y��I��|f=�I2A.lH��W�� \Y�(�-�o��_"l��hϹB+��������j�U�$�JH�\@dãy0:�i�hdJ8�W����]k��?#������v��jW���BT� h��_w��&d�8�\w�]+2^�C���~�vp�*{��y7��̑E,�EG��\��4Rl-��j0�W � ��V	��"F����}���E�~� ���#VJ��_Fu^DGZ���4W��K���3���6�c����]�y�~H�m;2h�N���C{��Ue��	��W��Oc^�z��9��Zv\�y�t��g�>:ɾ�
v_�.-9���������J��(�Q��������R@��f��701��J��/��a���ɛ��I�����p��A<_qng;��믖%�=�]}����N�s�/�5G@#o�객��5��P	׏yq�"�N�/�R�uv|�K�R9E��X?���ee���v�h=
��:�enh �fT4�Kn�0�{-B!��`o|Q����`�������V왹h�mcV�DJذ\��чU�[��������"pi�]�1#�iFb_�d��;1�\�� F/�x��
;�&}_��e�d|�xi-8w��O� �{�0�zι�|�u�xV��Z]�
_��ĳ�"��!�
��/aS�Bص+��H����_-�l+�m�h��S9���8�G]كZ��2n E���!�CIS���z�˷:uo]�CףE�b��d�Љ4��8���S�����.�;SH%�Ġ���Z��ҩ/L�5 5�c�8%��<�c:�m�O Jww^}{�&�ϑ,
�$�쾙rN��7@��f�����3s