XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>��� ��ZP
橱P�dB4�LI�3���A,F����%.�w��o��ڸF�TK��{��@�Ɔ�=<�����7]@`�lG�ȟ)Cw�9vV���!���yy	?7RM "���J�
�Ya'�(���9�ҽN@���5jt�Y'�w��]Q�����q�`&�k�#y#�V�K�
 t����<u���-!�ò�?Hw�q+|]�E�ξ��E�߃8/uW[[i�w�&cE3��]�[���	��A�N@l(E,[�:�����⦍p��h�[o��h���������۸�Rߏ���R����cܚq@�w7]�,O
�l8D���oϕ+c�W�?ɧf�|[�z�X�Ig_���`jn0O�V�ì;&�\ߪI��r��<�C�/~�J�@��t�m�ļ�N���ؙ�m#<|���qf���U	����R�pHea}����Pzr~(˼�9{cBK��/$`�"\����Ua�cW<#�!Ί�UQ.5r��y���V�Iߖ-E{61_xC��Jwm7����8?�t�O�w	!�Ĺ���=���;x��`�[}��f��b .m�lo��Ůw(h���֔��͊2��}�2�dJm-��Ϊ��A�+@D����jO��VF�7�ͮ9ج#�.m��F~�ǩ��rX��k��i�N�@���4?G����t���X���&���~�	��rk3��$���>���.���*�3�O#0У�9���u�
�:�L,ځK����������-�0@XlxVHYEB    4284    1110���PdɈ'��v���=�o(G�'��@=����2~���Hp%�S�ũ�Ÿ���$��X��g�+�&4�Z��I:-"v��	~k��)�z�LC��"����yl�)��i\^SV:(�V�I�1#@�
�^���hB��uH������K` ���r����"�s��nѐ����Ɣ(Ϥ+�g��;F�c,�
v��,�ِ]��40q�t*�4�-ܩ�c���\(��n*���!��3{�#��򽴾�mAa��}[���@�VtL��� ���xp��͐rB��b�,�D��ݼ��1�Z�UJ�{�o �ݢ��� ��I����>Dl��7���w���^��2�^N���K#�7nQ
#hA�W�����-���w�$z�=x�I*w9Fgq����۠�J����|7��{y
��>���~�柈n��!8;_K�������&�(s�o�5;2R�m<c���u3�bϾOqfl��5���GG5l���d�j�C����vP&�Ñ�y#�݁�Bp;���	��?��0���d��G�	�U�r~)�'�*���#���z�$����lg��&�Y'hm��W0B�cb�Mg1aF�h�O4��=[=ۅ�B���@"}& 4K,��<���ԟ��}�!,+8/
��<�5�9���_��7��2^׼?Eg�r���8�Q�ڠ>��h���y�Y���l��R:]"����R,]$ʼ��";,���Az�i�vƘB��'���T+$^#�=^��p�i��ۡ��/|������h��P�^Rs Ls��Rt|ˢ�^�`����������l	���f[�qOG�0����ؙ�V��W�Rs8b�dNV[���K�<Um9���*}�Ƞ�0�WMDO	d^�7�ʶ`�`h�*i��q���J`�A���2yW����u�h7���S|�,GFቧuHZ.&W}3�T��߬��!���\�R�F .���s��s�SSe�5���y��bY7J�~�ufm1܂\uAss�UV����X1:EÈ/������a\~��X*�[�@KQ(����R%��_5ܓ�)�	�Z�(h��g.�+z�x�}�K�G^�_��ד]/ɔQ�,�(�y�\�i��xa�ѻm��M�b
���TF�'k�M�ь�mh��.�w�̻.O� 25��E�
�L!��%��iL�c��"*'ɣ���N��!����	nU
C�Fǭb�`\���[�9TDV[���J+g���鰒*Ԃl2���i7Ą�l�{�v�G���ZI�x�q�̃|�֬@qό-� Y��ئ�퇴���&��@-'�GCHѕ��X�TS���P�J�}ʽ�"�KF�!1ɬ>��c9�
��b��E1���� �Ų�k0����|�����pp��i�P�C6�5D<��u^��_�(ˬ
6����� JTw�A:e�� �!,߸\��^���#�X�K���"�@ꂓN���������D�Kߍ�_X��~rVЖf�\-L�]A�!ͳH�`�\��0��P���W�g!M%Ѩ����ͽ�q�}��nU����< �g5p��&�*�Ԃ%�HQ���^���!{��],�[���cPI�aWA�^3��v��*;l@V4�q@��^�.FZ����u:���ey�k��f�:���������-�u�b��ny��_��3d_Z6w��J�%��[)�#G"�k��L����<���uE㥬^L��a	Ox���wR_e>J?�?oS�o¹Ļc�>j�C���Y1����&��[?�jmj� ����dw���&�W+�����݃���N���W���账{2}N��l��4K��i���F�GK2+��K��({�oۢ�+n�_ϑ����4L_��S��s+Y�8��p\F���Yk��c��r���^Rq*KFw7�bǎRh��<��B���j-j,!e+��0 en�e 0c����y4���h��v��SR�tb4Z����L�R��;6h�C>���M+ e:ƨ��}�{ZM�&��_
��2�k���F����d�1��W��!4B(�B[�mo�� $���c����5�����~�׃�y�Z�x�� � ��}3mǐ~W���2Sw��q\�z���׷�x������	��QP�����m	az���[��G��x�:��])��Ԥ7ؾTT�O�������k���>6���>ڀzS�D����ʘ�`lX�E��2�p�]:9Ѿ��)�4�st���9��#��p�c�:o�L����>�LX���!�0c��4�3���slΤ8�:�f$F�@�gZukx�g����P=g����pL�*&!�f+ ��*��Ei/�����{�`��f")X�^|!HL|)��[�fF����	F�Y���G���
���~@���N��e�%Y�j
�"oXܢc5ه��t�2ܔ��
�����H�V%BӶ��#�=�@eʖ������F.����{$7p�����*0���CW����M���ۦ�V6�H-q�ۯ��ƭ~y�&Ņ�F\��p��L^d�-<�$���vEfx�[�d�I?�Q�mۗW2=���	n!G��y�H��� ���H�;��b�D��>�w	$�m3�c�G�a�C�����ٿ�x�3�};:,b�,6��]X�uX9{���v�4Bn&�=p�$lUm���^��ݦ�D@�>x<��s|u������਎w��v�"��;ָ�b��1�#$J�5=�n���ݝ	0�P�������iy[o"L�h�V�`wP�����z�gP��30j�t�z���%h�C��)&�M�(7����������+�+G���.�0B�é�q5��'a��9��k[6`������=���Bra����Q��<��N]��0�g~�`���Q9��(��3I.k@��Z�|�}c@C��%ڄ�D�nkp��?�P���F*#-#À�I�h�sН���r ���N��}b<��l�!&���U�N�0Nb���"�H���G�^�/�E�8�����^g�$������tM�}\h���˝r3m�9�D��ht/oFba�J;㝁���<�����u�ۋ�[�)��d��%�Kpy��	�\�|�}��
�Si�aT�b��N��B��C�� �g�YKPiġau����z:*�`��U �X���Ph��D��5�*��fR�_Ƨ.�r�M�����I~6R[��3<b��d��5�10ט�����A�ٶנ��O��7P^bu;��EQ�^�K��ܗ-���*Q�uM?�^�W� +��0�[OSn���D{\��>�8��B{$O7ҍ�����A�#����w�謎Ѫ����b���f��^;c��Ԟ�ƛ ��m"	~�a�@�?j)D�W�L�͋��~�o��'k������N��7��,W�m��GU��У7��[e[/,���?�N'���7�;8�σS�N͘�3�ݶ���p����۾@�_9��YF�ͽ�Y2
��� �����n�ݕ��N���I��l�9�@U�M��d$�O������"����oh�"9"kjÚ�q�R3�SӶ�tH�� I�����n�k�pM�]dFQ���TНD�J`�r��u]�I���A�HT����Ҡ1蕬0;��KMv_� &j=U��cG���M���o�����r�SZ�h��= :d�X_��[	Xr��ua�sV���>B7x����O��5��j�=�J/P���d���l�d፻.���*Z!��_`������&�tB�gQ�C呍\d���rM�׎Yɏ�� )jAb��7~x����d���(�˞W�:��L���)]5D d����S�< d4ªC
��I���ґ`��j7��c�Mu��Z�ᝁ�60{W�zTtqԞ������5#��1s�+�ٶG̱}�Ce��������Cl���b���o ��f��	
�|:���.�3u���o5��i�K\��PY��bG�.��,Rh�3am����(7K�%�}6�J���dD�G2�Am(�6��-���h�UT,suc�=K�8bt��idTԀ��e� ����������v�'>O'%�([�<j~��8��{|�.�B3�ӣق��"���t��M����'%��O����f�[+T�8w��J�p���^�i��]/�L'C�FҚ�-:���JϜ�cWd�+�Ci�3��e���#�K�r��;S�	$ǻ��RH3����c���n&EU)�d�0�tkC�fXn
��b���M9,��,W��$Hy"8