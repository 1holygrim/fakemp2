XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���NR���!��[�6�m>������c!�3e���:��Њ�So����o�o�tXĈz�q�-��R��L_���g�E�CI=�"Y�j�θ�:�l)& |p��`Ʋ����?%$�C�pX�����B��͙���ATDl��\����Es<������t�Ykt�� �Dν��hI��Y��S�!hX~��K1(���|��%7��*LS���1��[�Vi&�)��l��c�$�$�X�%�惙W���H��|�;��U�R�e۴��N4��&@ٍ��3�GxTY�������~X�5��(,|K�D�nw&�l9�$v�t�\�P+T�3E����k�ⱼ���m����sʈ����2���eh��`��7����>ƀn����nZ!
9��d^�p�[�$�q}�@M��k2���-�?�U	v*�86�XcԈH ��3��Or�;��V#��j�M8�Q�0��|���҈��E��l�b�Q��Dx�U���P�͍��vH-QX�j�o�En�y 2�ϡ�g �w�7�K�`NM)��=�\ EH)��$1@�}ӗL�1!�0Z��ٮ��;�qO�M���-d�D��=oM�����*B��%�\OŇ���|YH����-��-~U4[�
�+����\̣Qq뷦/_y�R)S�xGA"�`guuP��W�6)2�=T��=ȞK>���:۾���;���MAc�f�~ lx�����u*��/�!������%*�� �q��"�ߢ6XlxVHYEB    9fc7    1fd0��;憙ơ�`��	����hg�k� �I7�0��#��T�:ܶ��K�$谕�4 ��;ja�����B��iM4;�d.滮�`�9�o���5�=��^ƀ��St�ۥ�ώ�/�!^dHx썎�r�v�z:i�'�\�zۚKh��Ιi	m�e�u*�5z���z�KY�^����գD{=�����2>�PEf\�L
���qY�BT�;h;��Zē~�d�<��᠄0�
.��`��RZ�d��ިQ�u�X���sD)9ԩ�`_&'��uD�M�K
}x�:��vn͢��|	:��1q�	��i,��d{�N�<�6�LJݳ��X�w�b��蘝a�C
M#��bf|��ܦ��d��?���V�%l��fx��p&'�'7UED?U����@c�	�}Z:곹��T�@��?H>O=^��)7E�ݛ�ꍃ́i86A?z> [�/�-�P(��t�d�2�N�pη�8H��_�o���)�s�֞{ԉ���Zӌ�ٞ!(]��/I���
�Q$ny�[ф�yEפ�t�k7 �l��٦�VP`��{�������+�03�{Y�fnQt��X�����%����P���W|k�@�T�V����ӑ�7&�� 6RjS���`]b{k�s���CO�)-�5�Ha�rO?'��J-��*|�����NU����sɛ����$�.��w���)��r<��`Q�|���`m�#ig��.���+E�Ķ���ˆ}��h��3��e��n���&9�9Q_r̋�i#��s����X�@G����ߪ��@���&��� ��M�OV���u���c*V���;��c�;E/v��0\�<����"�oX�u�̿�GM�S���j;�~�n�|1�"y��l GBC��-/6/tx�}�i�/V���x����25���۴�jK��W&Q0�f�4Tg�|�i�_JݡF(������K_f�O���7�eG����_<���ң(��*��	Q[��^#d����.����B��0�w>X1������J��2��`�ԇe�U&�J&X�H${ճ,6b���2E"k�Gtt���I���1A3�xm
ɠ<�D�V�*��f�:Z�\˜������M�3;�ʈ|H��VtC�Ք̼m��sP��E'�Y�����Ж���0a+�6z�T�CU�;�����M�w�����y����Aj`�.<���z}�~���3��"m9��B��BF���eػ�Y=�ڳ��1���xd��g�@+��罽�z�(� ���+��dBR �.3����vP5����k�nO=�r�Q�N@��$&*/��v�f���Ƽ�!)��f�b���c��qF�sD��-�ɑ8�ۻ������D6���	�U8��5�:ކ��r���>����AP��J�� 7~S7�li7���:bS#{�p�=��7i��%a�W���2'�$ J�A$@�J�9���M�J$_��2�R/���p�] �}'�O؊Ძ ����+w�4
����)��X��9�<�eōJ���u�#ܝg��LsQ� �w�ljȲ _c`���Iݞ+�ɠ�`�l)b�����RѐH�R2�d8��|�\|NG�d����f�i>�6?s2�D�D؄����Kb�Im��U�m���K���ؘ�Tr�ş��o�@ހo:?:Z��D�- ��j��:��S$4w@�/"�*�4r�6^n�[ћ��m�կ-��#���8�;Z�rZ�_K���o~�P�M��A�/T�dt&:�z���I&�?�.�*j#7[ ��;��O�5Gv�G2o�T�L�Q���1~��=~]�V#>X��p�5�K�����?w��&�����'o�9"=W!�s�v�����j���)o^�X�-15yhE$����H��]5�5Nv"ч�{n嵩�u	
?��|��G�莏�z�
�s�O1B��<U�m�@`%���D/"9�~�.�Z[��>M"�y�<��B��3-��KF��Uo��/Z��3M�c����A�=	�Ԩϛ+��vBVg��c�&�U���]��?g���폡�P���l�:`6�R�-��ƈ9��n��� u/r�l�*�z^��\W�&��C�Y��'Ĩ�3S�+��������,����P��F�v�0a���V�G�Z����y�u�0)�O;w�|����dp�����0��WM7()K�p�kLODߡƗ˷?�7��dԓdy&��Tz%��e���֌�N������VKpy���T��U�W�n�����`�Ye�`3��(������0,DQg?�w�sD�] �G��?�+Ue������d�S֥�p��I���H-m�A��\V��g~<������A ��OgCh¶g`|����,S�����&=�_�~N^^i�������#�괯�=ƍxw$��h�',�!/�
'9�:�hq������٭&b-�cjJ��W�(�	��T����R(�y�(\{ �.vU����g�����כ��W/���w}��/bb����O=�I�c~��9lLua0�Y�D*sؑ0Lf�M�4������k=�%Z��y�|ɛ悢}��C��{�3��K�e�YkR!x�"[�1����A ��D����m�cL,��˸�wU��O������8�5��7��֛T�/m�zWm{T:Y��M�\zh�Ư5�y
�b��7u˵��"��t�X�&����-�D�*N���0�@+�Z)ʢ�pc%]�zfV�{m�+R�D�U�UL��=lτ}�`)��*�A/��L] <u�}���ڰ��M��.`��:��6_L/�VEm/_��0'�6Tぇ�����elK�Y��Y	��P�o�KTC�}��z�Qb[B��;�<�K�v? ��S�K�������Ne�RF���E�eJ<.�����p���՜��븹�� 8�բB��O@�2�6��+�7|�����T]>D���g����	h�ƛڜ���� 4S��*9����7�]̈�cļ<A$|�����K�����P�d�Ŀ�WE>3쒮�)�`�/��D���U��M�W,�* ���.�]���b��Q2-&يXZp�[���k����24���H�k�{�^�foi�P����}�P����ºܼ�%�sb���羅h>� n8�~5�xf�a6�ң��-A���)?��z�k�b�Xg�`���]��n/���p�+m�ӂ���L	y|�-���pk<��F0ʥ�ܾhѺ4j푇t<X_k�)�w�4�6�����l�+/���
�Z�z	z��܈:8ө���� ��?�~O�˼�$	Eņ3{#h4a��|'�2	�q$�[�� qk�����%ҕx�0p����<�[Ǿ�6�g_{ (`���%�0Z�����_-�v!r�P���	Ge*CԄ�
'����.- �^i�߬n;���y���U��r�s��L�s��zf\�YQ�g4�������kiZ��@"0n2t�Q6���k�[�x�8>2��?�����Ŭ ����Sȩ�����U�,���� A��OXF�m%8Ţ/+����Y��qe���o�r�#����q7�մ@�i0/��=��w?6e+��j��A��&s�M�Зw��7#�^��G&�����7��W�V��$� {��]���\��[)<�ȉ9%#{�88�ʱ�S� (hG��V~)29��=B\�2��F�܁E膖��	e2Vhb Bɲo�&N�pL6��,`Ԡ��=�8���e'f�x�\vNF��3�r'�T}Z5�M}M�lR�%������j�)��U��ا�C�gC���h�(Z3��by=#��؎�Y�a X�5ԧ	u�'�d=�7/W�%m��q��z���s��t�!V�����w/��fto1� EJ�\f�¶iL2���Ɓ���]�� �\6�\n�$���������`­��G(�o֬́�����<�k��tC���OX!>{D�3O����A',A��K�69p)�a�Y�P���{L�Dz�K��%�8yz���Խ�T�D���")���f��Ā5ybb�a�YܼK��x֊����$�����T�잀c)�5�����r�?'b�t�u߸�$]0���#���ا؀Ż3ڑ�ᗁ�aƒ'E?M����8�'GBZ���Ga\qĥ@�L��������
̦��fhs!5|��\Lw='K٬"��mM5�X��r�������Ӥ%�#��m���4�:�e���b=ߌv�+�).Qr�U�)���w��BMi��,]�@-C��� c��?:���k�6쥘J�'
o������I����\ap�z�� �sx�^�~�ǟ��^����
�j�
n	b�b�!��>
ɒf���{.U�7uj�S �� lt�1n󼨭�n:�f{|�����E�Z`��Mո#����$�=_�zvBq(XA�d��g%b�4�4Q�C�5|�w�alwPg�<xʥ����a��D���|�(Q�������"C&4�;�}�Gk��.��(���toIN���v\��\,V��V���X���(0,�2�G9k6�7��I�ee0O�Ԏ� ��яT��{�K�.:gQ���9�yG-7ٓ:�:(l��� {�!��1�-����� �9{�L���A��9 �lƖ	�-]�W\"H6�b����ZX����nF��ܼ���ׇ-
_�p���P��5�w�߷#�BR��A+w��EO�����E�ۉ���� G.�+T���p���Pg69�O-]�d/E�.Ƒ��{i�/�����=&g&kZ�w��(es�V�b�+�$��h�;�>U��ՠu	,�Gki�[lغ"S2������7�U��a�ϯ#�X�R'�;�����RʢBM����e,7����'�Y�,�O�����+$~z?4� :7��)���%$Jσ<6�}!�f�V	��xŻSԷ��G���Ńw�sX~�(,gs�ف<Ě�)�Ox�������S�!J	�!)0�������2�]�2�N�No ٛ�I#�%��$*%�c���Ql#o�gri}7�v\�Q�7��3�*�nl(�.[g�6^a@�I�iJ{���V�]{ބ����n7��^���,7���b� )���?Mlz��<���Խ*���	���5�cR9�snC��G������|e��� 4L��!��ע��,����k,�|y)���l�@z$n]	s�NkEp._ԭ�k���ݹ�� $d�`*;�C�J>���n��;QM�og7��B}\�n1���RK����(�Ø���T�>9JG�����,�ܼGބ����w�����ȹ}�^䖉w�2�A�V=Q��o����a~gV [NJ�L�Qm�D����*|T=7�5Q�ʻ	!ɭ%������M�<Bܬ��v���?�=jLN�Rj�THQ$��%���P 1�G��	��l�q`˩l�x�lP��U����idf�:|k��/���<0��rorIz݄�˼���x����"~��FsŒ?��9Q��7c��8��km$\�X�"� (dv\��j7��)�w�)�<�')�P�z�?��t
[�#記���"��
A�#.� ė��J�E���#5�������*���&F��f�=g�WY��5�9����[j8
�����S�������@���c �a=�ƐFJ7�����P�:�x)8�i���?n���w��)��	\���+��&*�ؔ:����-��0���E����P� �������_C!���W��}�h���Ȍ�S4h�Zf��ٶ�h����˅�<,*�d��ѻʡ�D�w�q�AReb�	��jY`��q���	m=`(�K�J�L&�[�g��s���6��\�����Z��5��1E:���B��g�jl��(�w���X�����S��@��f�ظ���<�+�5d���~�-x�:�챌6��;j\*-�?��aYx`��X�p�-�R��5�1ε�[�&;r�h�\pqm���"v(M�*��X4b��J����"�/���Y?{5��0��S�d�b@k��j��Z)�^��M�0(l5jʽ�K���n�ml����諨F9��M��d���9d�O"�~-�ӢSV�db������Fx��c�T�t����e�ł�
����ԕTy�ޭ��N�E�;_���҄�)���kT��7��j�z�vXh���gKGVRYmW<|���r�~��R0j��$O���%�~�Qك��Օ2r��i����{!$4���fⳂ˺2��v����N�`".m��$ 0D���3�Y��U���v����қ�?ZN5[yط�Uf����i/B>� i�+qz� �Ӭ`[����"&���b�tO�?���^S4�Kk���pп��v6��.�!��O�	N�a���7J��M�q"4�ո��mv��'2��cčo"�����5i�ަ ��*H�,�`�LF���+�v<�$
�<6;������tX� �����4kL�)�i$)ܼ9B��N�H�T��Z:.�qp���c5���ǜ��S����<~��%&������dQ`������ա��~������+	{�< <1���|r���`62�:M�f�/�R:5�RH��'˂�r�_?JqB�X�s�N֠�r�$3�Q��D���+�h��;��us�L�|��}���}���d�˦�k�. ���,���P-5H�c�V%��a����yq�ط�YT��([I�zro1Ŭ͵�eC��L,���ޖ`�!yq���+e�1I\��&����k��>����I��>Cֱ��xD��q�$P��tXޏVZ׭�6!���=��n��5\L���~B�Ɩ����� ��J��;�S�Ϭ���C�n{,�d�4��W��B�)L�Ĺ�h��
,�װ��w���L�^úz^�Ea�'���7G�e�g��i�G�P���Jټt@ㇻ:q ��ͻ�Z�-��Gڐ*:��@���t:DGȤV?\�P�~�`�\*#9l{�{G E��\y�R����1��z>6�J?�*�)�a~�����-��L��ڻy�w׼��R��)�}C��Z��7���l����qv`���N��|x$X�̛���vu,���|���-�T�Pԉ	K�q��ՁR��#LD9G�ѵ��倦�	����]їݮɚ�?�Xv�L =.cR�� !(�WEN52,ָ��{� ���K�A��;V*br���M�Քb�3Vb�%)0����u�Gگ��/!p�e��0���ήet�^�@h>�WN�G�q,��14 �"c�����z^��rk����Ͷ�.P�����\v�����w=�"��|��7���T�jU���Q�s���,*ЉЈ��԰|䃷kg��u�p��$��U�O����)�c�
�w��G/�����H�E��ˍm�-��.A~�,A�G�kG6j}fML��Z�ɶu�9�e"b��c����t�ne���g7]W������+�4oAJkP�B�e�+��4	�1��������r{��i!}CZ5lH�W4�~־, S?�Ld#��F��CSP�?%�ܜ�o�����1�����n%t��>S-�s�4)J�'}�c��2X�S�G����{��׹� ���Ilbۤ��o�;R��wR����h�������w<Z)j�A��~˗� �+/������SS&���O����E�}!s�U�ki��e�S�\������%Љ���(۬Ô�Os8�>*��rRn�o�b�����s�[���*�6��,���J�AI�ZDF���{E�<��}��f��.���r��L\�������A�h��,A�s�i����x��2�������= a�������V��H��5���I�L���j}	}��'�hyV��N�譃d���l,��΀:8���?"�!��lmE@pn�>�"�ELo�J��H#�{���It�Rv���ֵ��Ő�$��6kR>����H���E�������&p|Y�o^	$��$�M�E