XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���������1(�1�5�4B���i�,�~��G��! �v�0R7�J!��������nn��kuiw%�2.c}�f��)&/6o3#m��W
2�=���v��9{��_� `f�������	%fXV/T�ZT͘@@��{��82:�A��.NG����L7򫂝��{�y���@/�T��5�r�E9��zb�MZ/p�Ց�B����0���*"x��8����0�g����"��7O����C�Q��d�)�0{�Yy�������,���������3߮:�-O5V(m
��J���|�R��bYJ���ʐ2fǶ.��z�g�4���d�����*���	��3bAjL�;8�L�w�������s��*�~�a���cuGp��7]��� ��������`����ۑ�$��_��������e�&���i��%�����H���#�n2��	���~���%��]�չd�mfc�	�����J�a�>��Sg�bf�LO��\z�����������/��вU��H<#�@ \�nUXW����zո �q+�ue={Qd/׬�4̤W2����ed�![.K����e����h�I��	�ԃk0��{�ğnCA!F� ve�.N؀y@���M�Q��w��'{�Ϙ1�Jɹ���[ ��AV���)d'P��?L�҅ދ��`�����Nʐ-\��Y���aKsk��^.j�GIrR<O�O���{�����)F9��k����`e��㱥�h�XlxVHYEB    b087    2540�Sg�74��LL���`����9A&��g�Q�z�J��{�a��<:�3Dq��%��p%��6j��z���0��eG镧��+�%
�ɸ�%f@K�>���;"*[}��"��Mf~n����x�.�H�p�/��ja-U���V�ٿ��>�1�]A�k�i��C�Xƣ�htG�5�F�h��ԅ�Fb�r8>1��=,Q66��{�u� �5f7����нY�,�l���,U����F�!��,��#>8�ٴ�� ¾(��?@��>QA�O��gD���+x,jI.E5�x%i�����VԺi��S�r�{��O�B�k�^�^�A�K�A��qT[E��4E�����c���Ɠ��4͡����$��<�\Gƿ��S�� |7р9��֐8|gbb�������~�O����r�7�3�'=��"勀\�y12�����x�z�0�d�:��+*.��U��QaG;�fmk�	��JT*�-a=e��J¤(�xF�����,G��j��'��B2���SJ�gy��9�c�9�E(%�v�C􊪎������[Ŋ<����#�ӷ��E���j�)�Q���'j��GW�)2����Td��3z�>UԦE��u��e�.裁nQtN����O������nVI R�K&�[#)��3�8ڒYvf�r��o+�z��{9��a����H@�n��Vv%b�1��k�wHs�]Ze�
����053��C�M�x�qꅮ�-�g�%m�K�����!7o �HF�!D�N%5���ߐ̉wl~o��!�@��7-�_�B�w&_�bN����f~Iǎ���^&9R�!!M��Jg��k�mB�>H�4'%�m��W,;�V�yYT��Y�<�V}��Ը*"���na٘����uL��y���6U�ʿpe��a�������ל(����bI�a���ꁆA���m#�w�;^G���� "d�Y��Pc�f�;~�"0S���%���6�=,�ƞ�L��C�����Q�D�����$̦_�
�1�~��^:��ja�%Y��8)����1HX"�ɐ-�;���٤ʔ8î�Jܜ��x���0���d���6`tN��l��߹h"0���oJV� �[!�=y=o�K|�y�.�P�ɑ�!�r�-v�����G?;�#��Yr�A�3�j���LR�rhF$���[wY�ֶ89VWҔ}������t|����_#5˲o�+
�E��O� �vF#�^��J1w���ݷ�a�B����ZZa,?3��� ��/�T�\l-�� ���0і�q|�A_j7'`o6j�yWvE��3�%MeJ ����{�H�b+f���²��WY��O����\��,�I�&}j�,�t�=��;E΄�g=r��Y���q�ƒ_ ����Q�2I�=慄v�/G���D ������U�S�V$�h� �%�W&�v$Ӭ�:��k�a ��{mIA�7��Jq�a7�#�s#������z<��*��c��mNgyt�N�z��&F���Q�8t>R+�9(�tڭ�{7�� �;g�$�=v�M4��]G����z��`�TBo���'5�K��SN���\�@G�[$&Ī�i:���%Ko�uW���$t�p�Ť�^Jĉ	r��n ��m�[D�4>2��A�F�Q$X�`�*��1����m
i�U��9[���T$2r�4�D��"X��Fg��)�'���q�v�yzN*�-z'O������P$�����Kͦw�	�T��nQ�u�+�C��櫌�`��D���Y���BF��:)b�gP��(��|j�%�
O�M6ғI����ἴ��@����TLiCI3�'�4��]�
e������I�4�ǃR��E����K�S����F����ڜ��簍�*�3�1Q��v����v�5P�$��!~7�Z����q���Y�a޼�:y��B�A��
]��D81���CP#��X�E\^x|g8����l|��E�;�@Al_ki��A�},�R��C���R�2���"N���
�1���V�n@�HQ�?2�%��<5���v�d[:�l�3aC���̩�r��Ap���2Vm`����t��ޡPŨQ0��(�დN�����I*��WS{y��W��h5�tדYN�C`.K�/��$E��!����z��*<�f�'�-�aEaF����3a�b�N�a��9�������[��#�1m���-� I����%��`��x&�iG��~*�y �Xb=*3'���)������=ƒ?暟.>	oO֟.��@վG7�j�#����cp�j�7U�hG�zT~6�쬘����V1��y9n�%�I;8_o��2�N�fT���c�+t7�����9K0��}�\jQ��23�~xڞ@��⯰*��$\����r����R�o?��{,^B���,ꆕ=�u��U>�3����)���i��v9�Ϧ�"�n��fR������(����3��]j-��1�)mF��W= o�(�"���5j��}�ˬ�����ǳy2�_O���	����(\�C��<����Ϣ��Y������;���pn�q2�@���c^�^����!�_t�y7~��R
KI�
�#�8��M�"���{m�^�r�2�jإ@r��d|��9k��x�3��c�wX��	pfMT\'suí~3
FF�k�����|�=�,(+nT-!��9ZVǵ�pk�
 
Bk�[K��(t��D!Fy��QĽĖ�厍�DUgq�OXRLV�J��O(�	VH�=E��$�)I��j���c/��/+�cT-2�N}�����Yb-q�S�5S>��}�m��Xy4[W�� �Y\a=]�����t�� �U8��y0��o=�*>�I��- ��m����GDs� ��?8��ZY%��]@glT��&�7�'�d�`7�SI7��M���V�~$!2���M�٘�t���TQ�6��+�cb\I�U�ctp�Q�Cݪޖ91���@��(X]k����n��@s#(K�/�8���"ˤ�L�r�yL��h#�JÑ�?:v�1[JgA�@)ʡZ��CTһ�Yr�ɃFtQ��M�\�y6�+�jf����J���&(p���r��EzA�G�����(.���
�k�d�z��"F Y�jS�����J��2_(>5T��h��,���Q��Y4��B~��Q�_y����@�ղv�E=t����	��D�	%�g�6�u�LO�(��-�@�ԟ�|�AV��i|�]�I����S߶|Z��ڣ�&�`d��i*�'H��:�d�9L}�)��褈i��L���Ǝ0@��ET���$i�;ê�<[�$�0go���B��Yw�FJ�BSZ�Ҡ����d��RP7�\���=�.�r12U�}`:�a9���

�8�C�Be%~��`�EndM1�ّ�qI�)}{����oS�-2����������������\Wū����QՙFŭ�j.>7&]Ka��[�)���B��:�	��D�'��q����R���P;��U�Lfњ�C���Z0�0o��6�mډP��1�[�u�m�:��Fd�T�/	%=�E%]ƽU6��(;ri=Ӱ����ړ����(��a��(���W�fD�o�������ʝ8��p���]�XR/��C�pqb`ͧi��T�k��Q���|�#�T��3}Y9��g�������Y�F�Ma"v]�o��A8�a��;ߜMnHF�úr�=F�@G�a��T�
�@� ���ښ���m�u�or}ż�-�kc�0@�K�VBF"��{랕HQ�~�˰wt]~cm ��2#I��K�`PQ��l��sGN���BZE��5�ރS\E���WPF�
��[u��F�rE�b�)r����Mk��!�[�pZ|���JK�t��{���$ԁŻa�>t]���,��/ȩ��$�����|oib����4X���C���s�=*�j���H��1<Ig����V+[�r�;�R6����t#]�uޚm�N)!�	ĸ�hnZb���9��J��	w���e�l8�g�h�&�K��#V�din�S+TO6�OvO�`+��zs&Dg �ܧ�˾��#Q��������kw[���*��U^��"Q\�g޼#>I���V{����T5��1ݝ���%�}�1�*!����Ew��5�Ӱ��|_#4����'fi�Ӿa���g�:^"�Uo�s�[�n}���դq�>�������׃(�)�GB�/���&%�����S}�HX(�a�� _\�k����}���
���hw}\�]������L��]H�=���2^��R��K5�	��G6r~���؇��/å�*� ��x�bG�A{Y�e�a>�����Swϯ�j��Jv�.�
�W�o�1HL^��uA��T��'�E�q-x��zk�H�iH��J�wm�"����OI�����
 OTH-�Kt���[Z�'��b9��&����h�����HL^���IX��m^� @�Z�G�A��W��� ��\J���'8�@6|ދug,f�܊A����q��Ү���n���E��?�yٜ��(��!��|�ū��"3�y^�9(4���7@�Ma5���<:*V�1N���;��S�~��ӤE*�0:��o��-W__��_�8�5rr��������A�Pj�N�}`�+*��o8HXaY���4C����j�ֱ�Dh#�̵���tpGmΠ�*Qo[HñC��Y`�%�n����_��hX`�#�>��BD4�p�Ӄ>�6l)R@2!	�&{E�L����Z�aಘ����K?��]�����N���z�Ssj_�mR��\k�n5�g'	S ���U!�@�	4P��L��N;�	�`�%�'�����:E7f�x���0�/)c�Dwy�W:)��b$4 I���ӷQ�*m��-$o�t]���/1D=㉣�
���<�AW�L�SB]�c���	EwZ�W
�k����2T��Y:����Q�T��/��7,i����x�W�h������l���Y�c��v-������%��/JsEڤRӰ��5z Uk�Áb��K\p7�q����\���f!ʏ&��+A����P��&:��v~3�d�9��N:��|��7:
{X���ì��4�XvcX��|HI��xW��"��(qf�,��6b��#IzTg��w�9MWd��S/(.ڤ�X�Quyb��-����Q�R3C��煱�U�pǠ��|�+�K�	�Ajۤ���l�
íK$mQ3�Y*�K��i@Z⣸憖��cs��Wz[e�h#����-8g�N��O��즽''��>���u^�(;V�������A�F�|��ၸCF�8�qHXrq���i�4'�}lߊ�1�_x &��&4��� ����D�ٮ����pۯ�{�0O�aXIh�w��u�b�t�|��}��Bf��G����O/�.��XTSG͍��'ʨ�6z�����g�YBf����p�Aw�
G�B��f�������U.�̺��UM���u��e`|��TI�*ҡ��=�4܆!������Rj�����跦 ��]�A��f�ұ��k�O�'(�؁��d�QӐ�x��	"5�h'�M�o��ްwC{	%ua`�D�8	�6X|2�Q� ����:�Ci5���i�o:������	�NB��J0(�]|<k���em]��������_:P-�s���t�ԭ t�e��jǬx9�>w�*��~��a��n��=V�u���_���5��c! �U_�~�CG�Nwy^ŝ�����0���EX�Xj�h%[�<0e��a�׎��a�7�
w~��# �AhSh�  �A��s^I��
r�?�25+f�2�a.Z��U�����$G�?Y��Zg���*�=F���q��z�7\�ɰ�Y��/�6��)�/3��K�����}��,��B_�j�v 1q���,��(�����=�]C &rz�(����Q!v���MtGF�d��FLiu5��Q���� ��+�.��E�v�գ�PKr�Sⵦ���"S�~ۿ�F�U���8%/;,a1cx��� �p_�x�M�sQ�jKm\��_�s+�.!8�q�x�pIASN��^�C�-.3����M6��z���O9IE��mE�F��ҏl�z����NC0���O �^��u�Ėǖ�^#7h��c6��;�߃����K��K W��_�+�A�Tx���i�?��6#���J��3b��{1P�m�ҁ���Z(�3B֏Ӧ9
]�?��W7��/���,��Z��?����9g�n�é��F�N	�DGP,�n7F�IL�(z���3~@��"��<p���+�_
�@���m��rd�� D����B�q�����j
�ގ��#�Ǯ)��Y+	ᇁ�V])��V���UI�(�!\�]1�g&��N� �P�:��`���3`��˽Q�JX"�ܟ�\~X�����,��G��}3$�����7r�׋���G�����Ef&��>��-���1���<x���;�U���C�V�⧐k<��������/�.(���ֳz���Y�4�iտ`(��5����^gy�
����/m៤���b���,a,��ѣ�{Dr����
�1�+3yG��s��U�,|���F5RG�A�2$�c�|�
��j+o�>�G�zC�N+��wr<�/�߰���u؀�ȥ �p�}�5~�n]��}�"+���Qd���/""����|��=VO��ɮ��+;������t)�����X����:�26m��~��iS�&�E�<I�]�<��K�pc�Uh�dugǏG&���MG�!?�%���ň�J�noÿ�$��7���Fwh��7�+�0ҕ%�QaEV��Vs��{�@X�r��B{h�&aα]�g�d�����9h���ˉI}=6�8�f@N�O��~Ţ�D|�K�ҍc�!�;�p@d�S1���и���q�%�֙л��+�g9�D��15��<���^�r=��:��/ ���f�'�;�k"@�	+��y��Ra�J�7b�?"�>^�NY�\9�$�>�O�w��'?X���8@$����
������}�[���ќ��������`M����J^��Q���nR�!~�m�Q�����x%��Drg<u0���<�uyG�@H���x�*���^�b+U�a`ۢ��JQ�?Lq�Ui� x�2��3TN���U���ξda]����VPp0�������J6�%ׅۤ�)����4�&@��.$Yp{����e�/�G��@E.��6L@����e����ng��H���ҩ{����@x\�+���\wQ	�f�� k��-�i�0�� �ʁ!Ϣ��B��%�B#	j�}���k�MZ��CSz]�N4��tj!pd�1�L���O�����3��{/�j�}lK�A�%-60oZ�[6~�:..$�8�|U��v�,���_F�E�
Lh��`��Z=2ǵ� h�{��/fݞN���g*�����u���0X[E��W�H������
���5����+S�:X���i�� y��U�Z������H�@��Q	�( �.�
��,���$����� i��W��^�͙Y;�4aۜ����Q���R4��S�{��_dڄ��?��F��v�p��x,!y/y�Wke�>~��^L,�Y��)�{��F�
k�h��fOs�����,=�"{F��������(�НA|�Y�[g���wGWg�+mL>�s��/R�Hj^Q~�(���h�
�?����?��w��'���y��hQ�0v}����d��@X[I�`�#�x�'�^3�U	���Ղ��Aȋ����
ᑂ�Oy�ѽ��ɞ�u%��>�P���8�R�у)=���?o^LHߝ644|**m�+�]*bA����E�Զ�Y�sx��5qG�|��*�o��vȞX�fl��ѿ�r1��^�zJ?g<�>U�x�7������\�qgy>�ښp�4]|A;�g��C��������p�G\�}!8�ĳ2���zÙOwK�诧���A�#X�t��"�E��#��Ҍ��Q,�Wg�QFd������H>��
g�m� N��w�l���Կ�_5��-���I�y��@K����d�֥
^�xi#S���\��(ʾ�׋:�}C<��׶������~��w*3+�f�%e|��̦ �l�2#�&�ͤ�� 5��YU�6�	ӓ9F8�Ihd�IRn�~y?���5'e(��m:���nbh��N�9�M����Xrf4N#�6�����m�@�љ t�3g����b�-��>������S���$�>�;�V���Iq���T,�Ec5N��x����f��Q��+h�(x��G(�/�<`�+��}�eG��J:�Q�Ğ���$�i9}L$�ʤ��s���7l*DB�Uhx;`�1c�;3�⁸���&�G�H��6�	'sw5��|�׋@$���5k��׋�i"��x�+�_a�D�Ȏ^���b�os�Ͱ�B�/��d�珷�|h��E���I���\:��~���k���"wfJ�v�_A���|=o�g{��?gz���y���G�pCj ��1z��Ó�A��3K�pz|>��Y��D�/˧���)�,��Z�x��(�pF8��?���D��Ac�f�T])G\���`�ģ�}�]��C��a�o�Zh��dTٺM��q�e9<1
���8УkO���5bo��G"\9��'���������|�Oz�N�W;)�D�>��E���]$a�H�-�k0��[O��/���m��;���c?��dnCҖ�#
c�P��$�SŻ�	�h��#R;���TY6�.Q���O���z�7���A�� @�z�B�=;��ǛX�)3�Z\
_a���Se��W�hs�H�M�P�-�ɽo<��,�V�* eً���ߋ����G��@������P�u/R�\��˹�����;jA�0�������ۯYg��U2���s�!��q"����� ���	�[��.>q���!�g����V���ȵ-"�[z�6Ӓ���Tm$�<��ݎlN}�J���cd�e,�NT~���f�؊�p[���za�-�}�ZkZMt�IP<&�@&5����w���
��
@W�u�&�,��Q�N�L����X��z�R'��9�d4X��${l�yC�'�KC����]�����|�1�`�V��Ŋ����T�Qn6gyS;xa���"����~@;3,1F���� �%CCe<)���u{�+���O:�[����_�Fޔ��|��z���%��l���mZV��B��gJd�
�Ϯ ѻ�j��d~*Hf�LV=JG�1���ɢ�{�,��\gr��,��&B)�+�\paY02�������֕w�M_��	:V~