XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������H�>� ��(��w���K���\�
�,(�p�M`��V��y�6�L���h�C6v�h"�1�D��z�V��7��* B(�!<�f���^:w���DЮ�!�Ȝ C) ���\cy.U)�ɵ\��:>\ ��ƥ6 \���
s��F�^��ÙZ��+E��`���<sמ%�{���?��[�� �lOU��Ʈ���Y��1�4� ��Pe����# ��$&mT��d��px[!����r�|�N���W�BH0���09�M�+�fU�	j'N�C���e��[�M⊳�_�ڊ�����:�Y��"b����\a�q�6?2iӣ�<�<A����ڽ�1�k@��nZ��?/U�N��% �]�V�6a��V�N�Hu$��T�����=ǽ��L�t��_����UK�:�+j�O뱹?y�5���A�IէWQ���L�5��+���v��~z7A$h�����&w��wG�+�ˊt�M���<-��l�Z���L�/� Y�s�(�R���T[��U;,!g�m���\*;�;����b�M ?� �4Ë��R�
@��_-$(of00Z�tݑ���;����BGVgfIK�d�ґR�������h�]�?���:�)�^@�Ӓ`�Xe�8�Ѓ�vs�����y���J�Ռ[uw2�rh�e�;�D��(�j�O��@욛wU �7��W�
O��z��t�r6:퇺�A�-RE������u,D��m���CO <�Dǰ��r�+̳���l��F���/*XlxVHYEB    da59    2e30��U�A��*���p1s־�)Ū�b��`y9MW�%�%��Xl��#Л�I ��=y�C�ց�*��y��M04 g]r�)6�*��^��c�WGψ��t��U�
��ER⛉\b{Wޭ�MR{kJpcKI���殇2��w�;/�Vk�r͜v�b�T��Hz��6	n��9,�	��	������TB��������q�M�Pp�{�Z-���s{�͍��b)1��tL��D�-�/�-m�{�5�\��4ȋԺ�y�E8}o�8G
v��y�I/�ЈdE��jL�ӭ!P�{-�?i��@�x.�L��<�<e��;����J��7���xH%�|�Ɨ��T�*���[����'�`?<��e��!_�H!��#/�!BU؀b����4H�~O�آ�Af��F�)� �k5��X�Fq�b��!f�����(����qg�qO�,����6��l��j���49+rP2`p3K`MW�A�ϊ��V>��9��\8]����L۸5�۩/X4{'밿x�_�i�Ŕ��҅�x_����Q�k:�b�}H��T�8C�����N
�z$-s���y�O�|4j�oB=�=$�Q�
���un�Mc{\DM�ºO�M�K�h�)����L.��9Ua��v�_\@�f��cA�Ɩu��R_*���e"4�%����h��W��53�E �&S�e*�#Ni���wP�X� &>�	y�^
�O%-5rxzN���Y���7��t��\l���CF?EK8�v��P�o�r�7�<R�*�g�X*��5�t�x�w��ܚv�f\��yV��UՊ��H�A!��6�<��2�E�`2<�P�[K_�f�ѐ�n��/���pӏD>����������������gq�<�����(�p@$�<�tѴ���q*���h�ӓxG�Uə~�\-�`3o�\�e������!6q���N���<3�g�O�$=GEy��GT��
�e�V�ϛ/��;��"��^��9@�V���Ly��Nf��q�2��`��}��͵fQ��'��N� h�R3d�ifs���n{>R@�(������F��wR@��6�5m���E&~�E���X��[zy��{wݴ����Ɗ�^��Jsk&'��^�58�>ˋi�ZG��d�Ia
K��k��R�Q�����5�O�i��8�ǥg������a&��s�R�a!7�jcu����1gm�\��<?yV/�
:L3C��@|s�)+["��J� ��_׎8��C�؆cUP\�)	�}���
���1`�Bh���C�ī�)�K����L�N�r!4N���#�i9������C� �����]��VR��Q\�
J��`\����M�9KN
ʛV�����7^*<��Y%������ �몄5sS�൬)d���T\��g�#M�M�$8ı��fo ��B>��DB����-�5^��G�kl�4�m�����n��-��9��40�)W<���$�[���RЂ�9�o	/x�,������U �z������z�z��t��"s�0��*Y�X��[�o�n��آK�i��Jx���u{��~<g��|SdD8�X"k���]l��k��g�K�ԓL�te%\�1{ ����׆��"��Դq$�)4��{��px;�Dh����d{�b�;�7s<�ו�~��>�؅>�RrX�3�]%����xx���V��!��K�>�K��0���'C�r䑳�N�eڅ#.a������/"�K�	Gt�&y�8��^a��cd�%�S�~{D[�u����ώ*ʃ�q	*�g��K�+���9Vk��a�*�2�"������㬕AC%h�mL�a�:����`��%�c�D�"�0�E��������L��6@´շb�<$"��ͯ ��öY�/���/��K���9)8�^~^J`�]���;>�����>Q]����]���fW�$�W����6ZH�Qhޔ{]��PGl�&A�ݭ7��\iR�1�Ia�骮ֱ)l���[e�K��-w~��h�-V��<��07����+�V����n�7��+�OV �SX����w��C�&�":"�枅��6u7���j�"����K�!JZ�w,4�w���`�h1ғ����d)���Zt��&j�5�[�%�Klֺ�Q��\����{R�㳵��_�Wg�b�1~���F���` �%�W@�7�P>��M� ��F�w�e���_}R�Ξ,|0�ֹ�^"F�Q��phe�m�K@[��c߾�F���7GT<���z_�F|`H	W^fO��b���gneaG���i�U�yK���Q�N���G9�)�����4!ჼ����]�ј�^,̊�3|m�� ����a�ls�&�b���}�{~�gAtO�ٞ�= �;ު�����?��'�Z������%*j���G����܄�J�|�*S��~�RN�r��s�*�͠�zh&fU@�l�K5�)�\����
�tF��:�p���u�a~�VnYDV�BZ�6p0�����4�Z�M�o�7���Br�+�m�[��5<�X��4�#���6RͨC�2WQ
6�yU��e��bş�ǎ��C�+{˰��
��F�@�!�lGο��0*����:���ή(5����kV�3׼�Xh�x#���vXQ �Y�X���M,��mC��j2�����e�"��s��T��x<���u�?�� !ZrcJmኑ�D�v[p/�܃��HhWerܡ�!3p�"�g��sxP��mF�Imn?�e�}P6� -*:���3Iq�M�,����<n	ɓC 4���|��Z���m~-�3�4�H�G>@�����q�9�3�v�(JQg�*���j�2�5�mG��<k�Fl������
����Mwy�8�!:F��Q5����8���|q���]�45uu8�i�~û�lF���น�x��)���8���� '�9�݁��Y�ecZ�(!�N�w�$�yE
�x'��J�����i[fx�ST��2t�(�o�e%���_52���巘F^���Y�G���º�c9�C�T��=�G��!2[qۤ�j���Y���ލ3Q��W'�J������.����k��z'��&�$�_�b��k#�Y�I�Xc?�%��rI�Z�e7�c�d`�|�uerI��r�=�����)T	��J�σ)D��A$�s`� 않1�&���`�n0����n�X��慪����͹7F��0��^W^�>MQ{yyX�	b�kl�@�	����eI�F�A{� �Q��2u���o�5g�#l��jq5��WҨ�w楯���qQ)BKZ��p@� ���|�D���lMi@�p-�J/p@0��=H�/�x�fQ�f�DZ{A`�{�g�����vs�<F��R_�m��c]w�2pv�tʡQ>Ж�L���@�ZW�<���� ۥ��8��	�E�B`�Em����xw��f������S_��L��`Auy�`؏�F��m/�/��L���Z��0%bd8S`w�S�G%�!������}7�Cx��=�V�QR],RN��p(*�[@��݆A�p�;�ǧ�Q��C���W��l���}��T��4����]����>.-\���K�j��.WlA��tz�ǣ�b���<�{>��W�W�TKEG�,�9�E��� �M�SV����Vgr �A�6aR���V�g����K�:�3;>V���w�V�mg@��Ѝ�7T��/��:��*,�}o�8g��$p�`�r�d>�k�(^}lMͭ������D^KÄ>b�=v��Ҽ�K�����8N��A��!�g��Kq)��'�2͸���v��1"b���x�*��������of=߱]��p�����9?YW���)� �!��`�s��{$����� ]]ː���']J3�r4M��p[��6E�^�G�i��W��;|����^�W�$$Vp�b�Q @ڟ�KZ��nm�����wZ+�ñ��k��J��{�(����=ԕ@u���AN5*h��@��i�������{�{��)�A�7>��?��If8`�u��R(�Rь���i�*
ݛ��.�å]�;$7Q#Xedû��$8���te�=	E��ĳc#���
2r��P7ۑ�^�'Ma�� 8��͗�*������C��Z/���G�Ԣz�T2O΁ށ�����86���L���"P�ǳD��"������*v��j��.�]!{�.�OF5��6u�DI� ��#���^����FL��0���8GB��p�"s�.r��c>Z�tҀ1k¨��H3����%�(AkWQd�:��j=;LxQ�cvqe��x�\��2u�T���yv�j���f2�����=Y9J�e�9�2�+x�,�{0\��G��T�&6j*^i�r���	�[i�Mf<�s~y+8���zG�= qj�j���uP9� [ԮS���E����X���5���<)8k��n�\~$e��9h~W�ÊS�^��m�V�*j�Xΰ�d!.1���o;�%���g�0��x�U��挠V9����8�?�%��
��<����c+� ���܎��Up?nSKУ�/}�P}mS�y-�N�r��Y<E@�Í؞�,��o:詯)�Y}z���[�� �oy�x}��ɶ�ԔÃ*���B��m�1y�D2�a���o���S<�qB��GU�E�v*��
��K��S�����*�O���`�P�i��i���B�r��U��P��>�p�(T�>�j��w�o�u~��; �U�]��֘E�3�8�4��~�z���� +�:�'߫X�UnX}M��Nd	�dJ���
���
`�G�vc�{<@���wH�;i�:vA13�|2�j/�����F�E�=,��-:��5��gC��q���5j�F����a�.���;�0Q���k�ҍ=�ΠiqZ^߄!�*ğq����/�sl?3�W��S�������R����U����@��RRJ�ݕ�r"�R�KH���DeV �W�*��n'h�Mx0!���8q9�r�g�-��?�!Y�E��X1�^�|�`������L��<US�v�c�vx�$Ø���Q��6��U��C&k����˞�⠿R�3zM:aY{P�J���� �ɡ��4(�%9Ii�&�Z��>)2hU/A�I���4��� �/ڠ�xϐ����l�.C�5Q�kXiy0������
�d��m�4a�R�=\tH�ztWJxE���p����8,?�4H�����Mf�c8d=Ob:�F0�ؒQUY(���M>�³����9ʳo֕A�N�3��@�2�r�V��8�v�d.t�DI�r�8�Y����g�o�b5?��)Z�w2�$�[�A.����	���+!G����>/���4j1>e�Z_2���� @n��\����>��M4����F���}QL�WF 3��5�a���*g@s�4��bHM�PM���&��U�~^q�6c3*�<Ӟ��O�&*����n���u�w�o�/9p���z�J�Q12f�aih��)�,W	�6w�!��į��Q3�C�F��	�1��yB̍�F��`�۬�%�uCŶ� �}w�<�0���J]ޜ��Z ����v�E�]@k�:m�^<��E�}Pe౨m�̹���D��R��-��(��;���DQ��dM�J٪R�x4����������o�_����<>���9�e�2�t��yvñU,!ĉȨ����Cy�`�0k�<āZma��lF��ļX������Y����<U�����G�{M,i�O�j`�v�vO��%g���+�א"��p����sS0���z�$�8'�R��ɏ<WԦh"w�c���j�*9(�g ��C���*=�un��!wT�Ew^`�]2�X�:��T�ų6�:'��	hZ
JT䋜�
�S�v-M�|C�g���|�g�p��0�`�qrd,�B5kT�1��;�煢��m{�O�����P���v�����U�=W��3�7��썜u����X X���=�-�0U����H.P��H�����e��,H��8{ې�aP?~��,�sXPe������_��1z9��Ī�<�˫�դ���h���8p�g����l(�/��y��1�W�{�"Q�r�������X�O�|N#�m)� �g��3�x�-s�:i�եбϊ�Z�Q�x��t	�S"��R+Rt2�P�������j)�Ix�Oީ�{Q�T��v!��|h���=�=O��H��2ƃ���["�Ϸ
���Ft���l��|)��dFu>-�P�M��1�F����JӒ��$���m=qN�&����ثB�+�y>�B�IK�EXo�4�eJ��$����*�a7k� %l���|~���9,�o5*~k�q�<�PJc�
N�[Σ����iIPT*���R�mn��ڇ%���l���z�8r�T�!JwZ�}�����֫#��jq�����'Uc<����(��m�~�;����S�צ��I�Y�������pc 	T�9��͵l��Hu/�T �|}?�q��4�2���*���sA	G�r���M���}S7�R�]U�?y��{�Q��ҺL��,kqב�~�yT@�ƹ�s��N�G��1|����2�Q�t�2�8CP���{�@U��طO�[���kE��b����t����O��Z�x&�i���[@�kl���'ҽ͈��}6�QsA�JR$7��٭M^L���?(���O�F���^��ΰ��8�ϕ/��mQ�����VD�d���Ј�%�ꔲ��$=���(���\�(q�k*���xE-ѕC�s�5��\=G�7�kGn&P�ZC�'ZU>����O-z�X�bTS����BI������-x���t�o�T@O�lK�$�������`	;�I�)��P�F�1�S���.X]+�(]<w�b�����U��s9�pJ4 �[32�̢�e��1��+���nK�����4O4�'����՗���A�w��H��7$.��E�F��}n�I�?���H�͹%�b�s1�v�)��T�8`�p����~���$[�r/�T��{�`�u�U=ަ��5��}cc��m>�c�b�5!t�[gn�� 4�|3���i�[F��eK�4�X�a}GxTN4u��`�M'i�G�S���/�]"]�`��a�5< �7P�c
�a�n:hѭƾ�P}�����B�Iި,��9��.͢��4'7�0��1M�D;H&��su����2H�Q�p��u�,L9�Y�r��=szR���gAv�Ж��Z�p ��4ȣ���e� y���/C�g�Q�&�\+[	6� �c�ka����sKN!;�mT�<�X�c�+��g�x�3v�YC�N���OR8�!w�`�g�Y�6&\��1�2��2���N��tt��b�|}�P�QG��iz�V���tW2H�!�F?hn��_7}F�B*\:��Έ+)���K�ʞ�aV��qi��Z�4��̰;�+��=+�*�Eƴ�N���9�Ի���H�x yxT@lwy�K�⅑\��0��"y���>^~>3d��q1���Q������F>?uv1�w�ޗ����ǟy�l��<���!����n��8�Y�L8���?R�T^8|�zO3й���VW˃���y�Ic���k����tX�����U�̻��`0�?�|��:�R�����Ji��-����*���ZHzρ�4�
*�{��=Ю�U	�� q*Ι���X�$�OdlVɍ�20�-�+�嬜V!��$�=M
�<x��Hܧ1�����d&�ص�Q[IW�U�Re]W:,�x�t��	��;0��% .���ԫ6n��:�yo��U+/hy��S�6���{�Ȫ��e�(���_��;1@���/���S9vD�?9�Y�	A3I�/wf�����bI�c���Jc�[���%���|'�-�W��iH��g�;�\'���bd�'��I0L�u�R��n�����z��l�>�#�ڌ\t�5T�]�G�͋�*AP�(���3���P �26�G��W�x�zRsV2�[�R��7%��U^�XΝ˯��)�J�%�Iwk�)�/��|}����N`6~�mhi��A��;~=7����"�de���>ZPw������@��	����Z(��u�)N
*w[�5� ^	=��t�B�������1�P�!��Z�ݔ�x��)��t)Q�K�^i����盌D����E��60���'��:��o�Y�$��+�K�)΍���e!���_C!�~��Aм����]s�d�)���׀n�����?͘�����/im'��0z�ql��?ʬ^'�0l�S���	\	��4�>��Hu}A�AKg�;(���ھ�����\�7�98��dsz5��)�s�^T,`��`�2�d�ÿd9O��8��1�n�O8б��m�to�c�F�eT���Yỏ�cR@U@��1HM2�@$Hp�Öd����]7h#i2 �KZ�(@��T��߈�r�� ��gP�z��UW�,^��ى?�� �e�3��ϭd�h��Lr��FP��59��=A��f�^�kX������zPw
C����<�|߈& �"�kv�"���?r0��8mNErU.��c8���I�i'ilȍX]
��$X����U׀��ʙ`p敂�������e��S�o/1@��k�'�`�z6�K���v � ��q�1��Z%sν�(�����l�)=?�~��{Q�E�-OGŋ�*��|[H*��TD# XH��v��`�
�cd�l� z��Y57p��^�`�r$$�N<a���$G&����\`��V�韑3� ��"�������i^������W4p-+R�;�U�D?��2 �50ۄ*�RUS��YO`Oy����
�L��L6���gs6����:��&�#7q4	Z��1'�/��@�Ј?��d(}��Z�9�p��\�;FWEm�Gı�4K%��QL�;&65*�F���i��j+�y��JH��o���4u�hxj�h�&�6���r֚��w�(X�[�����$�jǳc�*�1�q2ԽX�ގ�KZ�����TÏ��o<�\in� �	�w���������i��SX_�W3��҄"%�lɳ�~�@ۮ��2��d-���
���͵5�/��9��	�q\�kw���"ve"#�"y΃��F
�$md�܆��ɣFY1\Al�$ P��c~��x�q��f�b+��w&�/���Z�B���f
Wf㝜<VGp���:�O��u��kf���;۳��p+6��ҏE�k��}x���p�I��W8��RO�����o�
��ki�Mv%�b
�i�D7�l�^"�+��6�&�9$1H�_y�r����4L�S��=Z�_P,��2C\��.(���F.^��� 2J��w�yUPQ�p �]a$�{pC�H�q-���d)ŏ�e 5���js��C�:�apϡ��0�h�%��%㞗5oW6�8��Mg��Q��I}k8�$ɛK�Q��}���rc{���m��L��?�Ux�~PG��GM�*������k��N��xE2�1��]GI��ץ��a��5d�\O]kL�e?e����'I�T�����|j�҈nM�� �Lc*� �xS�Ā�~�Ŀ�DJ9@�9g���ꓱ�h_��d�+�zK��J�a�� (�>�|�ׅ�ؽ���,��!a�:M�Ą2��҇��L&��sg��9#�eBT���r/��S�Ԇ�q1c�:����F��k����[o�E,%��u�&y�IV4��y�a����v� �$��yUxЄ��	 �����u.�{���Pw}��{�|k���1�7�.���Y��)
����]A���6�??�(�C��@o�1'������N<<�U�r�j$����><�z?�{d�H	K|m~�π��яok��t]ɋ�����N�\Ӛ*Ut�_�>I�����n�tI��rܘ%��&-����J�Q1ӿ 3�:��.��'�dh���۩��V�B�Ⱥt��raPZ�Mk�=p��F� ,L<�(禧|�a�[C�E�A��}[�m#��ϝ�����D~��gb@����W�vT�`�Q��;�@� �\@�j��dA�iY�O��1!���)��#\�ߔ�p�ِ�I�Ll�؋��X5�Nɿ�4��yG�(�UD-��a�rF��zj��$���~���޷i6l��nd j��4�/�K̀D��0���(2^ީω��
�'I�P�Y6$��?U6���tCLP��Z�W����e0?�-�Y�}Bc4��С�M	Dy���>�=xI��A��ti�̈.�q��n4Sg5N[��a��O��]�~�T	
Jn_K�$x%�}���D�~�%#%�<�,�����q��h�(}��P]�\q�@1k}��g�U�����4M'u�1��� rP΀�T �%Wej�<���}9b���ј2�&�{����Z���Y�r�\Q1`��y�
��3�� �3�=&�g��ֲ����bS/����]����EB����:�n!:��J֑ u���#�؃C�\�r��S��/W����"���z�X]�����K�
^9u���8**�y�">Hpbc��{�My�%ww\u��<�l���J�m��CRLI���+�,��Np�y�ό�� �{��1��CF��t!���|�]�ը�5)k��hR����80$���[F,i�����4U7���0Rp6���'`]�O<�%�X��4=�G�"ۣ�.��jm�+q�z��8�eK9#������Ot*�{�<q"�8�G�h>��L�X�om�G�*�{/9�}7�y�ܮ�����C�^6��z��=%o.;. �Ɯ��f&#Kh����U���,r�Δ	6Z���� @gi��k��Xw�f�%$E�o>�>�`�0>2�`@{,Ր�4xCW��FYJƬ�1�<{��s���x�H����,����P�����Sn���HzExy�%I%��^��%�4�?y>9����Lw��-:�d�=�̈1���'�G/��d��<���T���������� E���43B��Ȫ����0C�Wg��E��yڅ���͑M�*��YvR�?D��9qkh,`]������|��Z�_ڇU�'�&&ڀ����!����C'��pjFИfld��e$qYoX�Z�eA�#D��I?�o�d7��a����-�dh�����!��fՈ���>0p{���B*V鈸p�am���3����a�Y�;����o��	13���m�z{�?���~���.\���)��߫�˟��4��=�뀄D����-�Ԍܫ�	=0�w�sv3�/L����TbՁve�Ɗ|�ں�T{������U��܊�L'�~�)�a4c�B������z ������!��L�؝�+��n��U��.Yrtv9ym����uN��۸E)yI�[�f���ΚdȔ�~c�w�X����,}^,��Մ��}���ܖ��Qi���w,pX~8'�f�1���U%ο/���˱��(��k��c��I�#��E�>��P�/c��w�&���6xA�����<il�p�d'�[` [�&L�����_����Eb���Q���#e愚�%P�Az�E˭���;�TV�6|/�Y,�:zg�k�տL��