XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��g�[$�*. �?BY$1�xb�.ܱ9t��&�ɦU��?0H��[g? �u68ɼ�b�*������0.\��<��l�X�&nK\�'���۪E��� �߶�Yr��a��{�Z�P(��"�"�bW�q�0�P"���/���6Jg��/p0i�)�KH��=�%M�ȣi\�W�r"57}H!�^�4Cfä���gX��3s#�U���#�o�B�~�q��S($���_�7.S�O��@f�j��Ѻ̉��ˍ��/�"E\�����Ȍz���NS{y��j��:"��b�.C^4^;?�z��{��Rw�&�	���)�j�;�%6�6T��gN���Z!�<�a��� W������0��@���J��?�2�BI�,*|�1D�ءFb+��@7-�SWӟT�4լ�S�C��Y� ��@.��v� ����Jlۙ�lgm�a�:xH]��M��~�c��T*�r'*l���y5݈6Fߢ�*�e�� �yk2���Wo� ��Z��,p�Dk,�C7����e�7�Ӗ�z��F���*��]<7%'Qh�1\�k��M1_�ޡbf��.`��>]��و<�q�(e��<B<A��Mf3��xO�	���IG���V߿O�a���)x}-���<S�q�h�p�xqB&��l��:��aX�t�h���:"��A�`1��!�ơ�v���v����KK1���O��f*��^�d�j��7�SP&b��D�F�dm_���z\�W%2K�`8a>��'��Ra���
}��2�XlxVHYEB    dd8f    2160�x�_fZ��zsN�!q(����-�ꆤa|=�38rz��ǈ?;�k��T�d�].8ps��F 8�W�	�+�n���ε�F�8:�	O-�2��p�<�4vH�%�-u��1��.�h�:	���6��l�?�sM�O43~�i��S�5��q'sfK�ᗫG=��?^o(xB��oM�r\��S��,[�l��.ɱ���L���g�ьq��%�X0�SNq���X�a��4e)��8&�ߜn~xv�Q��J������ҁm��)���er#2s�/H�2a�LB���3�C3|MO0uN�)��b3͟�異��GL�y� �=�og��wj���Ϲd�;������DfTJ�*����[�eP�h��v�����S��
��#�EC|h�w����x�V�H�ڏ��<�y��~��!���q����<Qؐ9�\?�G*�v�鼅_��b���ޱ%HO(,��\x
�x�L�g�Y���Pk&��,�]�gT�J�՞:ց��U������C�P4[#��K4~ZM�ݱX�N~Bj+|ŃA��#	�������Y�*�/~�/�av-0�	�8�t��"�4;��G[��6�L�;؟�ȸdBMy��şm� $�@dY��� H �r7Jo!����{�ÝϵM2D�R�|����dJ=u��=���W[I�9�{�5|`�����:�5�v�;�mJ�Zv�n3(��$���#v�f&*�+o+���8�v�1e�g[H�b�"����[�p9�:���R�-C^y��.r?��%��.�ͮ,�'1�gFG��XCЬ��?�Oh���B/>k�-^�f]��wN���e=3y�ˍ�D&^�}�?/��ȁ+Zl���;�#�ЄGw�`[��ȯ\ߣ���q�,�`1A�)o�	�N��Mw����{�{�pӲ]δyZ��=�����}B���]'���g�v�)МA��L}e��)�C�<,t��c�6^�F��u9 ���yR��)'C�@�� �ܮXOAĹ�s%r�N��]��+9�2d`A�	N�j�����8�ۃ*��O����(�,"�p�/72w$��a(-��	�x[OY<�=,Y(X4Z�=�=��L9���z��m
V��77�w��I�k9��5��&|
�P�>����8H�O{_�}Wu��(i �l�)��h���9=-�铀�,7��#��W�H�'�Gʽ\%_��	G7J2Z��fDbR�<�����x��ܷ��Ó^Zqls���մ�h���r����"���!���p��j_3oZ�����	'�T������I�� W<��-������*zl� �?�c$H57�!o�Jܠ��jS}�)pS�����:)w���O�zG��C�CX9,cFH�}�)�k�Nڙ���թ��vP�󻝦ĉ��D�0!f���>�F���m5�m��W�)�f�V��>"c;6���7d]��z�
eӶUI�^Xf�%�D&�; q��.Oft!J5���e^�H��y ��^�ś����D��|G<H����,�Ycx��0�c�c���P����p�j���$;r���AC�Q� ~��@�]b�*zC���j\/���,䡞�L!g7��aɘ��VU�r�h5��7�=_�12=F��6`�t��+|��
KBC���G�W����5�ԉ�d�¶����F:��fE�EeX�%1��ȶ�nؾ����1�%���x�u��K��X
��A��dC�IT!� �����)�;�F��ض;�Bq�u";�Z[Ej�0ݤ����|	 �Dl�>'�a�3��|bv�+��A�2V.��T&�;2��^z��������:��J�_�=������I�3����(7*�Jbr��GۡЂ��آ����),7�*�A)$��q�h��-j��������֚���j��x+����ҚpW��S=���ݶy��>Z�$$����Јn�3��	��Y`�@��0c7̶���x���s�`7s�A�q��`|�cG��	<6�O�xl��,�E%P�R�,�5�l�V�����8�ۜ���\2�����ʴ+�}�g�Ij�%�(>b��[L�T��a��y���Q#=_�F��N��������]G�6�� ��6u��kMAw@I�t�>��dak��X�j:������OJ�#�[
���T'W{ %�?�&������LH�D��k�km'{=b�Z�J��U0�R6\WM	܍�V|�|�W�o;�$0���'�w/��@W$>-�;<7��$1��C�F�Pd#
:/��HI�3ݲ�1m��ɝ��_#{��j���� �t�a�-��U�7���D�����)�ř�cR�T;_�ў���@�'Q�P�gCz�4θm�a(��~���O ]'�G:+g�N4XUiH��TP�]wLXH<2�~�%7'���Ra����o$�S�x����G%I;�RĶ�Xm�	Z�({x��a�;~�+=�/�G��b^J�|���O��Ɍ̢��S�`��]�\��h
<��{EL��Je~Z�i��A�S�}��D)t���_�)��!�����Q�ޫ�����&d&ٞnO����>�����{at���� �񄽠{1`+-Xϖ[���� R�#y=L�M_?
Yŉ���V��d��݀��3H�}j��Q\W�|�q1�Ѵ��/%I���Db��]�%��[��Tr��]2�%�<(TU�Rȋ|	A���c�K���������?R9���J�+d����N�h��dp�d%�C���*x����
[����/ޔ��)L���j�[�VG��b�	g9L�ÕB�w�X�oK=ο)���T��	G�v�ul�K��R�o����T���D9��sYѿ�d�^[6I��e�w�\�������EuSo�N$�K	��qj��8�߷aK�n�.O�\�v�b<w�7�啶4y]�<�E�|�ikB*f��D�oe�T���X�wD!1�����g�
�NKl�9�S�˘E�l5t�pk
}i�J���Y�7 l����r�.��!�L;�3MG��x���X��?�KB@�0���O�S���d�#xY���oX�˗�L��Uĭ3n�X1�v���/>��q�v��M��KL��4,�G��4��=�g�ǆ1	�YAr����$H��~0��;u��d�ʒ�!KN�`;�sL/�`2�N�2�_��Xc�T�/������]L�!�O=3Վ:Ϡ�s��
���9�^?��w��\d���Z�;!��RG��z�6�N�!�����֩���b����I��]	���H���iWT��K+��4����Փ�H&	��t^�;�i>:ׄ@@�v�@_1��7�xXe�Ȇ��VrLW�u����Ŏ�c��c�{��s�;��<�&C�-�B��y���J��ښL��f&�^�� m�s�|�\J]���J�6!��Q�~��,ʻ!q|��X~�y�"�U�! ]���ׇ��\��X���Ĩ.�(1��H�����9��t���orփ�-�a�H�COg[��{�2���lP-9�<:Jjǽ��|z�jV�9�T���IR���Oޝ|x���<;ė#6�V�}��������T���xi� f�VͲ�=M��_,׭��Wk�đ7��&K�8��I8lI�ZYmm�Z ��@o�7�J���Kh�PW��]{1hپ�����0*9��U�����Ǳ��RN�I�����0��5���1l* z^t"�5���=�GT�(w�@t��f�*Q�Dp�)��n���YJ���qcV�:�h&0v<1@i�\V�l���@a�dtI��?�j6A���ap6F��F��8a�<=�BIN��$c����s���
�UͭqN�\ۆ��0#խ�(q����RG�n�Ao�2�t� ��:Zf[fA@���`&~��z�^�G��8l��R�K�1!�����A�(A�m�x��tk�CpB,��s	�-�����)�S��;O�����s��K��9q�T����.�І���o���׮��'@Ҫ���;�,�q��2�u��)��T�YS��뽑K~rL�Uo7w;b��^�����w[��z�
�87�i�n;ؽ�6%�6X��Q+*������M�l��]���7i����1�of��l�ƭ�.JS��s�v�p��nO�8�f��h����>�L�*��e��ŕK����u8��̃�0�`q<�I,Qb��Y�C��A�I��Q�6�b���L�����h��,�?յE`9@��y�5��=#�D���!�"fX��>�7�Ʀ<q|�G�)���Y#Kz���LR���=�/!j�U;�E�:�؇���"Om^
`G��Qrƌ�]�E������`<2��Z'�U�����]O�H��q/�h��nSh_̭�����Ad*mN2V��rj�w�I�ծ��͡��%��$x���A�c��QV�΅{^�ў������Z�|�0wV3���O��c
[c���`4WØ��ᮄ�A�5y�>Ǚ>�F��a	~+�c}ᜣ�B�9L�Kz
B�e�4B#�O �ta�\b���\�`��C���^$g����Q������:D�[y�F���WnntF,T8�f^�qz@n�Gj�u�2����'�A���U>�!�2�k�!û��Ɇ�0���� 5��$z �=P�G�~=���:�{	IZzIwv���I�Tv[��!v�vE_�����e}4,U�d˯?����w���}����K�J��~�^������jgO����xT��Q��TӀ��8�n���\uW@���]VO������ɒ��| Z�KFp��i��T�n��@^����1��U�h�ۻ�N|�>�DL�#F&U�d^��de �~�%4G�(��RD��[tmh�9>BW��0ݓ-2s���йN��C[:�Vk}���#���!U� "y�%���[����$�{F��L�8��P����wwO\����'�j�����ɟP򸒙��ڡm"X�6�="v�o ���o�[�|�˵�Bgar@y�;҃o�B�I×�Kr�-3D�ꙅ�������!cX���s=ՐC��+�PQGO���́�X�Sv�\�D�H'�Mz��+TGr��s'���w������ì&����pޗ�19F��r�;�_�8rf�1��N�ܛv�Δ�j�q�p��y�ۿ�S%�c�����|� �i����ی0�7c�_�_4nʩ�_e-�L���#x���p�jv�j�Mvi�\D�"�Ev]7i�6���RtM6��Lf�S4�r+:��tg�t}��!�d*�m<��@��ؓ�n�.E��A�w���U�X�QL�q��K�o�k��NR��Z��aC��C�f
0��G�fUu�2A�����,llm,����;�_Fś�>mj�@��P��tFY��_�1/�B�9��RϏl�.��:`���U���"���>J��x�0KanD�E�axɴ{�J�M� ";#J�xj��{�+��z�T���=L��1�^>�u��G���l۳�t#�K���T���g2���-�	҂D�b#�n�p�o7÷�
H/��h���<��D�c�����}���Ɂ3��Az�A�r)<��[<�IG�wi��^�ޯ�X0��Vb��DIGS���Oc{�<��g������h.�#<�9��N�z�V��Y��x,2�p�Y��u�L�G�����Z}�����QteQ�S�٦�%"qH��h, K��1�%��S�F���ؘ�J�(X"��
&^�7ܦA���L�_��~��5vAM������U���b��U�iVyL~�r��*!�L�ؘ���\m0���Jd�S܌x��*و�~�����31\�o}%��㺾ó��]�/k��%�}�����0�_�?w8D}�H[�����
�LkO��x`�C`x���4j����b���/���c�aY��g�F�����G#&���4<I� � ��a:+��r��߾�S�r+Sr���D��%���q���%!ޗ�X(���B!m������@n�S;Cy��U��Q!X����m �c�ĻO����}�{5�U���O$�I�$���o�C����oEJO?,�nuy2m~'��	��у��x�C�����p[-���� �zKV�Я��� ea�� ���M���n�t�&�����̋X�����g|v��,��r�d� 5�*(Ƌܬ�ou �<@-���`k�����wFyѕ��L�0_m�F��#1a#��U��}���k�5��|zbO�E=/���?�͕�{�`�����}��<���-'�Y��$L�?yZ�|vޑ��-Nf�	�7�i)1���^}��e*-�ռO���������PE�s61Z� �`��A�l_;q?ӄ�:L�>1�3���MY>�6-̵����%$ra^gO�B0���b'���U�$��t^�R^��c}��g����f�1;�-d��f4R�mi�D���Ę}w�e>dh���y5�v\꿽����~�����⥴̶cx���$�\j�I�2&U����շM4���:��\�Ǖ�u��ޓ̍�1��8���V5��dP���B�Z_��P���Z]f�(l�"�j�����2_<U����8��=-���f����3�ʚ�G�)�j 
���o� ��bEyVo�3uͤ"�wp�!	�z��;�Z�`���~�e�K�?s/J�E��R)ڨlT�{�B��k�6u뇯�@!���6RK��������?�EZ���@���z�P�#\p��!��&����^ȭ�x �l�n�����;�d�^n�{��?��I(-t�4��4��Q|D\ƣh���������a�^����.�Y�(� ��X��_;֭!Ы J��EK���R�8�|8So6V�Է�yz����;ҟ��+��!�������&�I<�QiK�R��mrɲ٢��5xFmڢ��׺$���qņ��^\���C��U��2���a'5��xyij���a�PFGd�FTR?���Aj��mB���)�Z��K^V��Wk�����kh�@'��������E���z6�D�=K��$�*a�o�i��A���=H�v��5��)�����*)�)���.p�%��aс��-��~���-�[?���
��L��~-U�NBB�ˡ��؄��P���L-�}Wo�^��(o���&{b���S�W�~����i�=����;}�i.���7Z�,��Uz8g?�u�H�¢�Ƅ���9�t.ڀ�6����$a=T;�^�z����G`�b��>�9�#�NG}
��]_7I�ϲ�Z�("��)O$�W'r���m�J��`��KAf�����~�JE�@�N�W �֞ۻKFjUn��|��9ྩ������i{�?LSE|m��6VM��D��{��Ms��S,8�M ����2��SE��0$��~�����p �{�$E�R���N&�^;�k������!-�ٱ%n(}�gvM�4В������af��Q���&,V�����G���+d��n�Z/�''����٢��Mћ���}w8vi*~��D�F)��U��bdH"b��/^~. W���a4�c�Y賉T����$J]wN�ץ=�:ۏ�Ų.���.$I�W��JR�΀S~:Z�}z�	'U�xA��X��wU2k����{�P�N�D�~V�{��^�)������H܉�q��	�;O�L�����D ���Rq�%m�:�a^�n��\T/��¸3w�d����쨬�����PJ�]���B�D�y� �µ�ʈ�ƽ�U�������s��כ�����sYO[��r+�ViV:X���}�`b���tETw�ؼ;ϼ�1��G�}�A;�2H�8�joh���.��K��U䥊�����iy�:۞U'��Ӫ�
)��[�	��<1�	��a���Z,���C��.{ߣwT�C�|ْ��oM�sʰ݋Џ��]'�]��x�/�U����G��8_�'l3yA��=?xH-ᆕ	��C��K_�x��
O�ԗ��H	��%�F���焑O[�e�^I0�M2J�:�G�N���e<������������WK�9J�dK�l��$�꧹�v���&��2��b�6��`�L1W�Ӏ-�����޾h��5�[��0b����7���`:A��S�\�(�U��$�����!&v�p���N+�Zk�?Ĉ��qg�yV��=i����L	��g�к[����s�J�Ծ���� �ּ��D"�tڢ�$��|q�镄~�Uh�W#iA:b06񴋠�e���45��E5�f�͆�C���b��خD5���=U$ݝ�� �A����&�����&`�g�³"爘����-|��Jnw��\�v�����#�