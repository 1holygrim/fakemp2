XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���|�W���g_�A��v^��ϋJ(G谈I[���#A���?���R��H�b�lmr���W��p��S/*Z)��֤?��Lc��bn�T\�%.��}4�%��x�-���w �(j����ݷĥki.	���'�o]��c�1J0泣��C�)�b���W�'*�2��S��&�a��@m�muX"Ft�X ��-�G��@��ny�X�J��I�7��}���`��MͰX'� d�ٰ�?�}�?���`I�I��W����_n��ŷ��h�MפeUC�ߙֲ��Z�C�o�i�N�] ̳ζ�D%eW��_5
7�S���qC]�k�׼w�d�c��[�*�5u��W�A@.�V�8��Ep9+_�j����L]>��o-j-G8�6��uN�Y��B���ˢ���C����p&�U�hӜ<�ն��>D�����DQ�{����`+�p{�~��#�|=ý�~�@P�Q�������7�&�i1���1�N��Џ��f��"���Z�&х�2v���Q���(0#�wvT���u9P	�"��k��_I�"qX?K��]��z��G)�Z��~�0�Gl���^��g��N6�#�~U�?'��K+�)@x�XŬ�/uu&M��������޼ڹ%@K9r�k�Hm���kϲ�8�ʃ�;�V�A����˵N�i�T�z��>,�Y��N��;o�Kx����ɀ�[l�T@�D��;�F��h�MB��`�伸M��:��;0�e=�)7!"�<�	qJXlxVHYEB    3b09     f80h���Q����܌I�P�'L��R��q�`�C-����b��%�{B��'�(M�j#�!q��qU�\S�3�]x{�����TF&{�Ir���s�h= �b�h�˸
&�0�)؃c{Os�^>m�"p��DdZ�X��a��g��C���|��f��J��T���5�OSpN��-vg�mNdu:Hv�P��,߶��C�:�A
:��1�Ӥ�.�F��%�[͝�9v��8���AM�e%������+��:����7�!��9u���>�<FU#h=�;OQ��g��#��#�E
v����w;��Y�o&Rj�AT��!�����C�(�4�
*����G�@q:8Ҳ4+n�	����}k#F��h^��SF��1�66A�R`������T�r���	�J�ޘ#
���t��SI��to�q�W�b�D�j�]�i�)��Y
����*ŉ�;�=����8��rj�v$���j��dBf��F�GRh�����J�� ����tO���󰛼�L�Ad��`���䜹����6\��/پ7�Z�.`�^|fW�AjhB��\�}A���);X��NSSɑ�bd��L?1��K3���ꚱF�![��*5�&��s�#�Mb���v���[x���{���s�Ў��C���P6��M���R�ݠ��-���=UT�Z�1�00�����*�#Cx�@���x�d
�J����"��BK�=�G�p���XΗ����<���'C��ӛaθ�� �Q/��� �8�E����G�@VU+HmȦK%g�]�@2;-��n�����זX�J�aق�/6�7�6\�`%V�=��FKg˩�L]i�VҦ��|6�>�ۖ��夒�J1��|5��IU?1�])�
�:�_��ͭ���9���K1}R�����2赬v��b�2>���	��D���������Y:�?��pu�I:a1�;�Β��^�J;]Iȭh�N����9�(c���_����:��R� Ѝ��<h�jmT8,�R��ׅ[�iUP�����-�����\�
�-�h~暊@�Ĺ�����|8C:v�Ut.>��=��͠m	�6o�z�/��X��Z�����x5l�U�((��i�f��G�:��]�C&�~��VN%X�� 7ȇ���/��Zj�9�)dM�+k"��.Z�C�T	9�Ӧ����i#� G�r��Cz�E������Y!�"u���_a�6�F�?��1 �Ĵ��	�Q� �r���?��BT�QA8p�	{�|26G�4�������S�UB�uv���SK�{Ô�����1}0
Of��AA��!a&�\����LuT���nn���5�S
����o��ݑ� T��!MY�_G��U�"�_h����PX4�Ӫ{KL̡�S��g�6�w�b!�q%�4�S���H���=���f@���?C��Yʟ��G%��V��d#7�NvhF}��ׁTk̆\ ��R��){i�ɓm���S}��h{�	 MPv��e�%s~�>=ov�c�����h��� �1��+�M�w�/�Z~�\�]�Vͪ��3R��_��b�N�6+M���g��rv	�%��
ou���k#*s/��b�9q�������ky�Q��5�&�ni�ѩ���Vֿ	�U�Q��94F��;�L	ߎ�p��q��v!�9��8cWK+1�y� �-����:6��X��̋s���>2����I`�$�Y�K�����-�+aYKbe������RZ���o��|�
<Y��).��c�U,6^�Ɋ�G���o�
jC�IK��\�N|���JK�r����P����(�%��$��R�m���3��\jY&�w[��[[LxUIx)��?)���8T��Q�"��`\.��,�A[M6�ŕ�<1��|<	%�C���1 a!<��m�Uo��I}27���ح 	
<��bԑ��E��a|�:�����c��Z�CS�C�Q����Xy73�:�x�-�':.f�S6昳��[���NK��Z\����"��I�XN\���x�Bx&gZ}��ۼ�r I�u��`
�ǆU�a�C�~@��8Y���81��l�����ؿ�1Y����9:ڕw�U��w�ވD!�G�P�q c�����k�6��/*|���.�ϻ��9��hR{k�Ã��,q�6�5�*�N�W�:&3nv�dw��f�ԣ\��;M�ʦ&����v�%��r�!<�������o���%��5FM�`��ʦ�r<�P:�/Z�phi�iU�j5+ϛ~8̰2E�&�}o�t�φ�srQ�:`�)����MI�����GN��R�#g�;�I��[��|����w��g��-L�8�6u��!�I?+!�{�;D� �{����s���p?F�q�HJ,�r>�&$��(���\D�XV�O���݌c�%����H�u�9�md|zT��h-+/��nJ����L�j#yh��)Ec���]�f+Bu�pY��!ϚIїg�a����{M	�Yc�����
�)<���t�(��*w��+%����KA��I�0�SF�̒��?ޕXa��1͛5*dH�M02M��m`֧���X���ȧ����¾�x���s�t!�T��������[�h�iG�  rI��v���'��*�V��Z���34�Z'S:�]xƆ�Q��+{�F�ڶW�"�Ry�E���@�=���A�`�Z���D��4�$��6d:R�I�L��i�ܿ���]K�V��AW7�O��k�N��Ir8�`�}o�p��9K˽��{�<Q��3��6��g�b�j�V�F.H��:4����o%1U7_�y��I1�;�Ҫ���CɝN'���F��bWlm�K'�n�M��>V	F�ڕU_�=��Ø;�BS6�=v'1�Mx�Zy�o$�G�9��F�/4� �,bL�����CQ*&E���{%^�Kl��*��ki�4*�k {�+&���!�^	��y���8�+�Wv�6�7wE�pzj�9�E6�8��l���*��J�75i&.�g�g�\-{�>�O8�YƶW/�3������!���>D��0ధG��#�e/Ƒ�Q;�־$�퉝�°X�C��|�4b��:}�{�!Q9k�.v����;�@5�1N�z�����U��$f����o�T�?�{8L����s>�����S��(��E�W\�>5w��؏�R�\@��)p_�w�d���ݜ��uT�2�0��A�R ��?��gS��  Py�0o����H ��:��'C�0�ڮg�T@�Y��ŞB:�w{Ɲ��k�$i݇�%Pg5�A�� ��=��R|�>��]�UQ��53�D~��w�-��+�/���S�ڽ����1�����|@!igGI��F�)�O=*��x�R[[�MC�l�� |�$���f�V���,}��l���D;S�U�nτ0�r�@�s\>y�?�[��(Ɠ�kg���ў�LNG٫��h�]*�;.�\�(qG�hJ^&A/(�X�����_�>�	��Ș)��ԋV0�(l�s�1��i�� ������=�Q� q�?~؅w�ؖ]�:�:"�
ŃY9Tp���Ǟ�x5�)�SYC��8<iЉ�!�|�d]�n;=[������BݪHz"�Z�-9</׵)5�֫��~{t���eЍ��+c-ra��2��89E�-W�@
��Ī�p ?�֓ <◢?��GO%��%����}����_�g���w{)*]����A�3�ceB�~�E���'��w��Ce�\�\Y}�u�wi�w�W�@Ol��[B֜�M�%� ���7@�l�lU&������^LF�l�7k��b�":�Ю�ʴ5��1��0&�h�oc��٪�)�L�u5j��ͱ�P�7���hUD�