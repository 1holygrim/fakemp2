XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����|L:I��y)>" �L(�t��;��e�w��	�7�T��siR������<�j��I�u���S�סY�8�)�9^N��1!�&�uں�^+�Ҽ��nd����ŞG$$|�h�M�)�����Z��؈���L�`a��C�K&���ߘ(�@�}�l����=75��[�v�̷��E�^�ى"�z����{��fA���4�h���sB��)��l��ٴ���H}M�N�0K}�7/8q���7WpA͸����z����k�sXUgYĲ����9w��UL޸x��G��x[��|�_��2�16 e�5�}�T�0B�M���m22�:�S�5��W��8�t-��d ����u�A=��SN�}Q�ˀ�Og����L�"N�*'�������v$��.8�a��&�!L��5�cȀj�n�d�f��fh���Y|se}�&V(@�SX��c�g݇ z�,�V�n���S��ДɎ�=�P��D���~�H��2��k�;L�د�k�C$�;X��*�d4��hJ1�׫K����5�Y��@�5um/[y:��vO6\l3�e�X��z~n�R�H�<RM�Ü]�`6(∬�,W��m�I�jvbp
�1� Qhw1��c������&<�s"��q�˧��a�OH��+>���%�x�~�.*b��?�T�$��3�I�WL�T�U�\����E�q�O�2mDA�+SUv4#N���|J�	���XlxVHYEB    5224    1740a0\ő�����c�C��1��-��w�g%�Ô��k]K��  (~�MrC��X� �w!�Go� ���S̞�g���N�v��g�
xF��n�������G��j�+}�UZ�f���T9�bj���7���wlAV㴑~~������>&��y���(x��yNd���sf�4_��EF�	l��3YA'�����wܾѹ�Ӗ��y�����vu=�e~�S��,�����ċ�y���v�6���xפ����Em�	?��`箬�;v��զ�X��r�{{P�LT�{�;Ժb��q�!�JLLIv�PY��N�ʃ�fO�gg>:�,	�CS{?Yda�O��-rn�J�k��mwac�o:��8eM�Vcp�|د�kӟ�.|V�h��%�-�1��yjg��R�p�5�}��b�JW�:,S|�w�ٯ,���v�߁��,M�h���M��E,tԏ}sZr�����KTc�H��k��eK�i�t�e+�|�M'K�l�N>!9�����E��@h�o�A+2�'�NH���Eq٬�G�&iw��3��C
��5Ɵ���/������c��yɯ�=�+Uy��ߵ������x��
wpu�ɛ�Vcٯ�(ܶ�ȉ�	\I���q��K��+����n<}���$���t��F�R�9��T�:ܶ�Zý9{ˆ�>�5�)�9��1TA�b�9:4���ހЂa��T���΂���f�u��=�$�G�gv)���e��I�u�weI2�Uzb�!�T�k�Paur������ok1*��gtoR)1O[�2�x������O���<~�A	����Ƅ�!h թ�	�g�Ef�(��!�Y�K��O[8�W[��_����
����-Ũ��W	1��?�T�7��!YJ���3>�Z�m����VDa,t�%r���z�~��i,�-w#��C����hq#Kj�n�J���Fye�:����+�0q��bFd	A�T�iYn<xN�hK�w�׈S�<�4*�ﭗ����o=-��q��#�����N��%<�D��i�k�����+��^B��@Ұ���-��T�,}/�m��aIe���I5C5�/"Yi�$�_�c�B�ҧ�=T�ⵋE�`�Z�Me��ξԂEj��E�>;(�������$�%D�&�oO�bf��y�L��8_���4'�
�t|f�J}+n��	�T�����҅+B2����p��2#9���=�B�q^0|E��i�Y��?I��Er�o�9�4e4I�T��L�)V�����@�����c	�vw����D�����jϜM��Rn�"�Ӭ���X��[��nAS���.��t5:�1qg���^g��E�F�a����hݘ2G�s��/)HS��lӼh\��` Z�_X���� >�R���n0_���Ӥn�t^�`�5w��~�D0a�[`5�^��R�֕���r����5P]�d��و�@�����Q��e|M&���(��m�x$�Ǖ����Ƅ��L4���75.�z����F`�[#��DQ�|]�����]�-8*4����ܼ1r5���e�y�q�QL��_D-����v��o�v��lV�o�$�AP�?��`#J�jF����R��ږ��s�:<�n�����Fڏ�	)M���Pº'�u>PN��U_.�3�D�M�3=��x��<�JH��[��]�P!h���I�E�m��!�b�+�����cј �<L� ���d�q4�؉O�����3(�Cd����A"#��~�{��K��{؀�u�?]�!3-o,6�{��o�MQ&���
� ��4�)� ���P_p�ɠ����i��e���w�r�y�8�#t�PlO�S��o$ ���x)��=��Q���(N���N����QO�N��܃�/�k 0�a_@�"DZͮq{ӵ���F��=��WE&��5�<�myvѹ]�!N�l��Z:�|�W0��ˌ�IA�i��AR�Ά�U�����
���BT(�q�������XSh�2e&D�c�&C�M�a��|�6;r�T�务�b�7w����vi�`\���`���yFFi�MY�i��Fm��d��_/7%<H���Z�z,�,��l'Q�	��'ː����q��IGj��K�I%��Ѥ��c��(2&/�>�`�7�t6֨M7<߄�+I����Ra�7��'b�Yg$%@|��f��s��ٛ-�|��b��>��[��cS�t�\kV��~O�O�q�,����[�ȯ��=rQZGy�8�X�a�i�\q-��	l|�6�D��i.1:�5���'UI���e�� �;���d(,�@�(Je�Ȫ��i�l�v=���#�U��1ñ<CH�5z��:�ǖ������ς_�i���愚,͕�a�"2�OR����Xo�"F�qIrA�!k�z�Ob��F�&��=�~!b�N;����=�	���l�au�s�LΗA��ۙ9(���}qc�:��z[��3������)�� >b�;��'�3uͦ�W�(t�|�C���zP�xʎM��;l�&!r�q5,�u$�S�qmD��ęS
��>A9w����z�]�;���PA���{ے�m�"��~�����J�1����/	>G���o^L��O�%9��3q�z~l�tׅBt�K6����bP�ۙ�F+�D_������K08�}��0���Tk���x��f0;�S8sU~���W� ��kf�h�씨v:�9yw��9+&|5��2J̜_H��6&`�\+�5�����t�Vaw��i���KX�2��W%cv��>HV}2%��#��aG�x�w�7�t�G̀��OC������-�Dfm��iIB9��0rIV��P��d�]�7�ǽ���<��f�=�|w6w�q)�Ֆz��^6�6<My�T�>��ˎ?�'�'c, ьn�zU��Z�Yu��Y��3ՙ�o>�d���"&����e�P\��7�)����)��Ý��U�I��I��7ת�Ll�[�dp�l�ߚזcF�G%���qPL����Z��U�9P7��+���n���T�o�9��G��#��z�ѿ��̰���"���X;�h�<�#�*C�Hímk�MQ��r?����B���F������x� {�(�v\hE�H^��2�(�~M����|q��<�J�\ �ε�Sp��w� ��F��@�b��]�B+jċK�7m$�#|��87@a(�c��-)h���ny�<r��R���a#gW�O"^pEC+�je�a�R}2�i�P���ԫ��8��0��$��p�d�9B#�?�ߜ�!�J�]^�@����íܔ�!u��br���E�7�����4�֤_MuA�E�r�&�4[���ĹYf�Z�����{Y콍�@�#�24�)�3�"=�6r9����Q�5�>3{�48%���nv)JA-΍�h��-b1(Pnoc����o�Y)�eT ����]�����]�����LF��\z�w�������T������+U�U� ���z��
�%5�R�"<�JZ�Ҩ��rn?��O!� )�dD���e����l��XYۑH�(>C	��DI
D��b�t��M�x�7��a����V֚����1=��coz��6*�10?�l�F�Q#J��o����[�2^��߸�@�ⳮϸ�xK��<�ߐQg;�������k2�|��C�;���rs��Ai���y����7�kY��0�]��w��)EQS�@��I�[�9KR�S	IGU�Ⓡ�jfCf�HIcك�#f$����Oc�t�]>eT��G�F���Ѓs*�-%V\��'D��,������1]M��!	e�B�=�D>���&zac��o�ބ{D8�I%'�W�G�4�1I�Q_������Z�!/�Ff!�k�.Q�����49���&�G��'˫���o��8L~��{���b� ��(6EA�X������B�q�E�9����z����ѳ��'�����[^��ps뉞�;��.\��u,Ľ��r��$Ў��^u�>��������=5�2i9L�,�@��Rل�1}��v��nM���E��b�b�r��>N�w��W��b�`v�����{�a�w��/���Ұ2p~�2N'�I�H��&�L��r��Oɕ��f�*j���9ۗ�����a�/@*������b} a��ra`?]���~,O�58Z�XD�l�o��2��j�ޘ�>M��R�8�=�|f��LL�>�=�0��Sβ��o��↎�����Xɬ���ܕ�9FlB�����=�6N�ͫ	5�p0q_^(	����|����YI�V�3˻��li�3�7����a8;˰�8�ߎx�8>��)<?����q1����m�^��P�qفQR���ԁ!)������ӊ/��f��GY�^��=;4:�1�P�&�\�Q����g�۳���B9M��{.�y�$.r/g� _DZ���d�u��
�x*j��a|E#�>V����q�4l��/G�=����Zv�&�]]��(K
~ �?S����+Cjj��=y�Y�)%�;�/��8[q�1V�14��6�,)*��L��>�Ru���bn\��|p�2�J�Xw>����aŷҼ��C- ]!��@��BW�oɺ�6��<�����Y�榎��&�	~dks��w���3�{��촘W�Z��&�a��!v�������S.۾q�E����P���F,�6�`�,��
D�4�Y���?\������-J7o��B�HPN� P�SI�Tw�����|��Å�'�r�,����7�t�(��f@����	#`���y���v��P/]���n��7�-׹�=����,�Y
e"L��/X��L��t���al �K�e7�%����u�X���ƶ��b'�q3"4Re�d'u��2n���֚B%�DB7�`�5���߅��T3����m���P�4���'D�뿢Uj;�m��Q����	*���4��D{9ŋ#5�'|&�E�g
� 
���t�XÛ��|-P�����k�SO��,���UXrJ�LU3/oU�iA���-+������"�?��w�7���BO�[�=졀�);�M1��*rQ]Dyԧya`g���ce�@�+{��U(%�qG�>�.�a��Jf�PR V��gG\w�	�C�A��hV�ݟO��!d}ȡ��Twq��[@c�H=�^����g�v�����g�]*��衪�߇�UvQ��A�y%Q����~�0Cm%d��c��HU_w��	&���K���Nn@>�U��݈$���^��<���3�P�ڈ�,y>�ٗ@�j޿��o]�-��[�\(ΐoxA7o���#3{a�M�XZͱ�֐�C���P�֒��E�P��lܝ@�[%"^����z'q-C�칤> �����APG?1��Q�l�R{@\5���&�ǧ�v5��Fe�M���8��Rx:�"8�,�l�&mS01y�{�J#0����?�KT 8r�&�M�O,C�b}�:��]����Ф�V`����9)�{��n��1'�X�R������"���µI�Ǽ����=�3A��L��Հ�������Ѩ��V~�9�J�q��Sn��_ؗrxQ�}\���'�zb(����#C=t��k���2��� �� Ar�_(��7�鮊;��|Kz�:�j�u��N���i��,��vE�K�װ��7��<"���P���Ǧvn\���z���h���F��νH�_'�7����n�,H�$� ���l-�o�-N.��$��ס��\�f����z�3]t�a���kɅ�x,��a�4�؄
y���m�583?	��c��h�����f�4�A/F�H4#3���f��o&E-�SL�E��Q3�(.��U�Y��f���z��Ӷ%K�B^�b��~��